module opicorv32_control (
    pcpi_int_wr,
    decoded_imm_uj,
    pcpi_int_rd,
    mem_rdata_word,
    decoded_rd,
    decoded_rs1,
    pcpi_int_wait,
    pcpi_int_ready,
    irq,
    decoded_rs2,
    decoded_imm,
    resetn,
    clk,
    instr,
    is,
    mem_done,
    next_pc,
    reg_op1,
    reg_op2,
    trap,
    mem_do_rinst,
    mem_do_wdata,
    mem_do_rdata,
    mem_wordsize,
    mem_do_prefetch,
    pcpi_valid,
    decoder_trigger,
    decoder_trigger_q,
    decoder_pseudo_trigger,
    eoi,
    ascii_state
);

    input pcpi_int_wr;
    input [31:0] decoded_imm_uj;
    input [31:0] pcpi_int_rd;
    input [31:0] mem_rdata_word;
    input [5:0] decoded_rd;
    input [5:0] decoded_rs1;
    input pcpi_int_wait;
    input pcpi_int_ready;
    input [31:0] irq;
    input [5:0] decoded_rs2;
    input [31:0] decoded_imm;
    input resetn;
    input clk;
    input [47:0] instr;
    input [14:0] is;
    input mem_done;
    output [31:0] next_pc;
    output [31:0] reg_op1;
    output [31:0] reg_op2;
    output trap;
    output mem_do_rinst;
    output mem_do_wdata;
    output mem_do_rdata;
    output [1:0] mem_wordsize;
    output mem_do_prefetch;
    output pcpi_valid;
    output decoder_trigger;
    output decoder_trigger_q;
    output decoder_pseudo_trigger;
    output [31:0] eoi;
    output [127:0] ascii_state;

    /* signal declarations */
    wire [127:0] _5442 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011101000111001001100001011100000010000000100000;
    wire [127:0] _5421 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110010101110100011000110110100000100000;
    wire [127:0] _5400 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001011111011100100111001100110001;
    wire [127:0] _5379 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001011111011100100111001100110010;
    wire [127:0] _5358 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011001010111100001100101011000110010000000100000;
    wire [127:0] _5337 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100110110100001101001011001100111010000100000;
    wire [127:0] _5316 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100110111010001101101011001010110110100100000;
    wire [127:0] _5295 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001101101011001010110110100100000;
    wire [127:0] _5275 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111001101111011011100110010100111111;
    wire _5296;
    wire [127:0] _5444;
    wire _5317;
    wire [127:0] _5445;
    wire _5338;
    wire [127:0] _5446;
    wire _5359;
    wire [127:0] _5447;
    wire _5380;
    wire [127:0] _5448;
    wire _5401;
    wire [127:0] _5449;
    wire _5422;
    wire [127:0] _5450;
    wire _5443;
    wire [127:0] ascii_state_0;
    wire [31:0] _2615 = 32'b00000000000000000000000000000000;
    wire [31:0] _2613 = 32'b00000000000000000000000000000000;
    wire [31:0] _3664;
    wire [31:0] _3665;
    wire [31:0] _5190;
    wire [31:0] _5191;
    wire [31:0] _5192;
    wire [31:0] _5193;
    wire [31:0] _3743 = 32'b00000000000000000000000000000000;
    wire [31:0] _5194;
    wire [31:0] _5195;
    wire [31:0] _5196;
    wire [31:0] _5197;
    wire [31:0] _5198;
    wire [31:0] _5199;
    wire _5200;
    wire [31:0] _5201;
    wire _5202;
    wire [31:0] _5203;
    wire [31:0] _2614;
    reg [31:0] _2616;
    wire _2619 = 1'b0;
    wire _2617 = 1'b0;
    wire _3872 = 1'b1;
    wire _5182;
    wire _5183;
    wire _3891 = 1'b1;
    wire _5184;
    wire _5185;
    wire _3947 = 1'b0;
    wire _5186;
    wire _5187;
    wire _5188;
    wire _5189;
    wire _2618;
    reg _2620;
    wire _2623 = 1'b0;
    wire _2621 = 1'b0;
    wire _2622;
    reg _2624;
    wire [1:0] _2639 = 2'b00;
    wire [1:0] _2637 = 2'b00;
    wire [1:0] _3677 = 2'b00;
    wire [1:0] _3882 = 2'b10;
    wire [1:0] _3880 = 2'b01;
    wire [1:0] _3884;
    wire [1:0] _3878 = 2'b00;
    wire _3881;
    wire _3883;
    wire _3885;
    wire [1:0] _3886;
    wire [1:0] _5143;
    wire [1:0] _5144;
    wire [1:0] _3927 = 2'b10;
    wire [1:0] _3923 = 2'b01;
    wire [1:0] _3931;
    wire [1:0] _3921 = 2'b00;
    wire _3924;
    wire _3925;
    wire _3926;
    wire _3928;
    wire _3929;
    wire _3930;
    wire _3932;
    wire [1:0] _3933;
    wire [1:0] _5145;
    wire [1:0] _5146;
    wire _5147;
    wire [1:0] _5148;
    wire _5149;
    wire [1:0] _5150;
    wire _5151;
    wire [1:0] _5152;
    wire [1:0] _2638;
    reg [1:0] _2640;
    wire _2655 = 1'b0;
    wire _2653 = 1'b0;
    wire _4132 = 1'b0;
    wire _5034;
    wire _5035;
    wire _2654;
    reg _2656;
    wire _3356 = 1'b0;
    wire _3354 = 1'b0;
    wire _3557 = 1'b1;
    wire _4758;
    wire _4759;
    wire _4760;
    wire _4761;
    wire _4762;
    wire _4763;
    wire _4764;
    wire _4765;
    wire _4766;
    wire _4767;
    wire _4768;
    wire _4769;
    wire _4770;
    wire _4771;
    wire _4772;
    wire _4773;
    wire _4774;
    wire _4775;
    wire _4776;
    wire _4777;
    wire _4778;
    wire _4779;
    wire _4780;
    wire _4781;
    wire _4782;
    wire _4783;
    wire _4784;
    wire _4785;
    wire _4786;
    wire _4787;
    wire _4788;
    wire _4789;
    wire _4790;
    wire _4791;
    wire _4792;
    wire _4793;
    wire _4794;
    wire _4795;
    wire _4796;
    wire _4797;
    wire _4798;
    wire _4799;
    wire _4800;
    wire _4801;
    wire _4802;
    wire _4803;
    wire _4804;
    wire _4805;
    wire _4806;
    wire _4807;
    wire _4808;
    wire _4809;
    wire _4810;
    wire _4811;
    wire _4812;
    wire _4813;
    wire _4814;
    wire _4815;
    wire _4816;
    wire _4817;
    wire _4818;
    wire _4819;
    wire _4820;
    wire _4821;
    wire _3660 = 1'b0;
    wire _4822;
    wire _4823;
    wire _4824;
    wire _4825;
    wire _4826;
    wire _3760 = 1'b1;
    wire _3752 = 1'b1;
    wire _3746 = 1'b1;
    wire _3740 = 1'b1;
    wire _3737 = 1'b1;
    wire _3700 = 1'b1;
    wire _4827;
    wire _4828;
    wire _4829;
    wire _4830;
    wire _4831;
    wire _4832;
    wire _4833;
    wire _4834;
    wire _4835;
    wire _4836;
    wire _3808 = 1'b1;
    wire _4837;
    wire _3871 = 1'b1;
    wire _3938 = 1'b1;
    wire _4838;
    wire _4839;
    wire _4840;
    wire _4841;
    wire _4842;
    wire _4843;
    wire _4844;
    wire _4845;
    wire _4846;
    wire _4847;
    wire [2:0] _2607 = 3'b000;
    wire [2:0] _2597 = 3'b000;
    wire [2:0] _5204;
    wire [2:0] _5205;
    wire [2:0] _5206;
    wire [2:0] _5207;
    wire [2:0] _5208;
    wire [2:0] _5209;
    wire [2:0] _5210;
    wire [2:0] _5211;
    wire [2:0] _5212;
    wire [2:0] _5213;
    wire [2:0] _5214;
    wire [2:0] _5215;
    wire [2:0] _5216;
    wire [2:0] _5217;
    wire [2:0] _5218;
    wire [2:0] _5219;
    wire [2:0] _5220;
    wire [2:0] _5221;
    wire [2:0] _5222;
    wire [2:0] _5223;
    wire [2:0] _5224;
    wire [2:0] _5225;
    wire [2:0] _5226;
    wire [2:0] _5227;
    wire [2:0] _2604 = 3'b001;
    wire [2:0] _5228;
    wire [2:0] _5229;
    wire [2:0] _5230;
    wire [2:0] _5231;
    wire [2:0] _5232;
    wire [2:0] _5233;
    wire [2:0] _5234;
    wire [2:0] _5235;
    wire [2:0] _5236;
    wire [2:0] _5237;
    wire [2:0] _5238;
    wire [2:0] _5239;
    wire _2635 = 1'b0;
    wire _2633 = 1'b0;
    wire _3945 = 1'b0;
    wire _3539;
    wire _3540;
    wire _3541;
    wire _3542;
    wire _3543;
    wire _5153;
    wire _5154;
    wire _5155;
    wire _3582;
    wire _3583;
    wire _3584;
    wire _3587;
    wire _3588;
    wire _3589;
    wire _3590;
    wire _3591;
    wire _3592;
    wire _3593;
    wire _3594;
    wire _3595;
    wire _3596;
    wire _3597;
    wire _3598;
    wire _3599;
    wire _3600;
    wire _3601;
    wire _3602;
    wire _3603;
    wire _3604;
    wire _3605;
    wire _3606;
    wire _3607;
    wire _3608;
    wire _3609;
    wire _3610;
    wire _3611;
    wire _3612;
    wire _3613;
    wire _3614;
    wire _3615;
    wire _3616;
    wire _3617;
    wire [31:0] _3585;
    wire [31:0] _3586;
    wire _3618;
    wire _3619;
    wire _3620;
    wire _3621;
    wire _3622;
    wire _3623;
    wire _3624;
    wire _3625;
    wire _3626;
    wire _3627;
    wire _3628;
    wire _3629;
    wire _3630;
    wire _3631;
    wire _3632;
    wire _3633;
    wire _3634;
    wire _3635;
    wire _3636;
    wire _3637;
    wire _3638;
    wire _3639;
    wire _3640;
    wire _3641;
    wire _3642;
    wire _3643;
    wire _3644;
    wire _3645;
    wire _3646;
    wire _3647;
    wire _3648;
    wire _3649;
    wire _3650;
    wire _2627 = 1'b0;
    wire _2625 = 1'b0;
    wire _3811 = 1'b0;
    wire _5170;
    wire _5171;
    wire _3873 = 1'b1;
    wire _3874;
    wire _3875;
    wire _5172;
    wire _5173;
    wire _3892 = 1'b1;
    wire _5174;
    wire _5175;
    wire _2651 = 1'b0;
    wire _2649 = 1'b0;
    wire _3941 = 1'b1;
    wire _3944 = 1'b0;
    wire _3554 = 1'b1;
    wire _5039;
    wire _5040;
    wire _5041;
    wire _5042;
    wire _5043;
    wire _5044;
    wire _5045;
    wire _5046;
    wire _5047;
    wire _5048;
    wire _5049;
    wire _5050;
    wire _5051;
    wire _5052;
    wire _5053;
    wire _5054;
    wire _5055;
    wire _5056;
    wire _5057;
    wire _5058;
    wire _5059;
    wire _5060;
    wire _5061;
    wire _5062;
    wire _5063;
    wire _5064;
    wire _5065;
    wire _5066;
    wire _5067;
    wire _5068;
    wire _5069;
    wire _5070;
    wire _5071;
    wire _5072;
    wire _5073;
    wire _5074;
    wire _5075;
    wire _5076;
    wire _5077;
    wire _5078;
    wire _5079;
    wire _5080;
    wire _5081;
    wire _5082;
    wire _5083;
    wire _5084;
    wire _5085;
    wire _5086;
    wire _5087;
    wire _5088;
    wire _5089;
    wire _5090;
    wire _5091;
    wire _5092;
    wire _5093;
    wire _5094;
    wire _5095;
    wire _5096;
    wire _5097;
    wire _5098;
    wire _5099;
    wire _5100;
    wire _5101;
    wire _5102;
    wire _3547 = 1'b1;
    wire _3544 = 1'b0;
    wire _5103;
    wire _3668 = 1'b1;
    wire _3678;
    wire _3679;
    wire _3680;
    wire _5036;
    wire _5037;
    wire _5038;
    wire _5104;
    wire _5105;
    wire _5106;
    wire _3787 = 1'b1;
    wire _5107;
    wire _5108;
    wire _5109;
    wire _3698 = 1'b1;
    wire _3692 = 1'b1;
    wire _3691;
    wire _5110;
    wire _3693;
    wire _5111;
    wire _5112;
    wire _5113;
    wire _5114;
    wire _5115;
    wire _5116;
    wire _5117;
    wire _5118;
    wire _5119;
    wire _5120;
    wire _5121;
    wire _5122;
    wire _5123;
    wire _3802 = 1'b1;
    wire _5124;
    wire _3794 = 1'b1;
    wire _3793;
    wire _5125;
    wire _3795;
    wire _5126;
    wire _5127;
    wire _5128;
    wire _5129;
    wire _5130;
    wire _5131;
    wire _5132;
    wire _5133;
    wire _5134;
    wire _5135;
    wire _5136;
    wire _5137;
    wire _3810 = 1'b1;
    wire _3277;
    wire _3274;
    wire _3275;
    wire _3283;
    wire [30:0] _3263;
    wire _3264;
    wire _3265;
    wire [31:0] _3266;
    wire [30:0] _3267;
    wire _3268;
    wire _3269;
    wire [31:0] _3270;
    wire _3271;
    wire _3272;
    wire _3260;
    wire _3261;
    wire _3281;
    wire _3285;
    wire [30:0] _3250;
    wire _3251;
    wire _3252;
    wire [31:0] _3253;
    wire [30:0] _3254;
    wire _3255;
    wire _3256;
    wire [31:0] _3257;
    wire _3258;
    wire [31:0] _2663 = 32'b00000000000000000000000000000000;
    wire [31:0] _2661 = 32'b00000000000000000000000000000000;
    wire [31:0] _4993;
    wire [31:0] _3756 = 32'b00000000000000000000000000000000;
    wire _3757;
    wire [31:0] _3758;
    wire [31:0] _3792 = 32'b00000000000000000000000000000000;
    wire [31:0] _4994;
    wire [31:0] _4995;
    wire [31:0] _4996;
    wire [31:0] _4997;
    wire [31:0] _4998;
    wire [31:0] _4999;
    wire [31:0] _5000;
    wire [31:0] _5001;
    wire [3:0] _3856 = 4'b0000;
    wire [27:0] _3857;
    wire [31:0] _3858;
    wire [27:0] _3850;
    wire [3:0] _3851 = 4'b0000;
    wire [31:0] _3852;
    wire [31:0] _3862;
    wire [27:0] _3841;
    wire _3842;
    wire [1:0] _3843;
    wire [3:0] _3844;
    wire [31:0] _3846;
    wire _3853;
    wire _3854;
    wire _3855;
    wire _3859;
    wire _3860;
    wire _3861;
    wire _3863;
    wire [31:0] _3864;
    wire _3829 = 1'b0;
    wire [30:0] _3830;
    wire [31:0] _3831;
    wire [30:0] _3823;
    wire _3824 = 1'b0;
    wire [31:0] _3825;
    wire [31:0] _3835;
    wire [30:0] _3817;
    wire _3818;
    wire [31:0] _3819;
    wire _3826;
    wire _3827;
    wire _3828;
    wire _3832;
    wire _3833;
    wire _3834;
    wire _3836;
    wire [31:0] _3837;
    wire [31:0] _5002;
    wire [4:0] _3869 = 5'b00000;
    wire [4:0] _3388 = 5'b00000;
    wire [4:0] _3386 = 5'b00000;
    wire [4:0] _3788;
    wire [4:0] _4547;
    wire [4:0] _4548;
    wire [4:0] _3696;
    wire [4:0] _3694;
    wire [4:0] _4549;
    wire [4:0] _4550;
    wire [4:0] _4551;
    wire [4:0] _4552;
    wire [4:0] _4553;
    wire [4:0] _4554;
    wire [4:0] _4555;
    wire [4:0] _4556;
    wire [4:0] _4557;
    wire [4:0] _4558;
    wire [4:0] _4559;
    wire [4:0] _4560;
    wire _3066;
    wire _3067;
    wire [31:0] _3069 = 32'b00000000000000000000000000000000;
    wire [31:0] _3068 = 32'b00000000000000000000000000000000;
    wire [31:0] _3673 = 32'b00000000000000000000000000000100;
    wire [31:0] _3674;
    wire [31:0] _4968;
    wire [31:0] _3672;
    wire [31:0] _4969;
    wire [31:0] _3371 = 32'b00000000000000000000000000000000;
    wire [31:0] _3555 = 32'b00000000000000000000000000000100;
    wire [31:0] _3556;
    wire _4670;
    wire _4671;
    wire _4672;
    wire _4673;
    wire _4674;
    wire _4675;
    wire _4676;
    wire _4677;
    wire _4678;
    wire _4679;
    wire _4680;
    wire _4681;
    wire _4682;
    wire _4683;
    wire _4684;
    wire _4685;
    wire _4686;
    wire _4687;
    wire _4688;
    wire _4689;
    wire _4690;
    wire _4691;
    wire _4692;
    wire _4693;
    wire _4694;
    wire _4695;
    wire _4696;
    wire _4697;
    wire _4698;
    wire _4699;
    wire _4700;
    wire _4701;
    wire _4702;
    wire _4703;
    wire _4704;
    wire _4705;
    wire _4706;
    wire _4707;
    wire _4708;
    wire _4709;
    wire _4710;
    wire _4711;
    wire _4712;
    wire _4713;
    wire _4714;
    wire _4715;
    wire _4716;
    wire _4717;
    wire _4718;
    wire _4719;
    wire _4720;
    wire _4721;
    wire _4722;
    wire _4723;
    wire _4724;
    wire _4725;
    wire _4726;
    wire _4727;
    wire _4728;
    wire _4729;
    wire _4730;
    wire _4731;
    wire _4732;
    wire [31:0] _4733;
    wire [31:0] _3546;
    wire [31:0] _3551 = 32'b00000000000000000000000000000100;
    wire [31:0] _3552;
    wire [31:0] _4734;
    wire [31:0] _3380 = 32'b00000000000000000000000000000000;
    wire [31:0] _3378 = 32'b00000000000000000000000000000000;
    wire [31:0] _3314;
    wire [31:0] _3312;
    wire [31:0] _3320;
    wire [30:0] _3308 = 31'b0000000000000000000000000000000;
    wire [31:0] _3310;
    wire [31:0] _3297;
    wire [31:0] _3318;
    wire [31:0] _3322;
    wire [31:0] _3293;
    wire [31:0] _2659 = 32'b00000000000000000000000000000000;
    wire [31:0] _2657 = 32'b00000000000000000000000000000000;
    wire [31:0] _5016;
    wire [31:0] _5017;
    wire [31:0] _3791 = 32'b00000000000000000000000000000000;
    wire [31:0] _5018;
    wire _3695;
    wire [31:0] _5019;
    wire _3697;
    wire [31:0] _5020;
    wire _3699;
    wire [31:0] _5021;
    wire [31:0] _5022;
    wire [31:0] _5023;
    wire [31:0] _5024;
    wire [31:0] _5025;
    wire [31:0] _5026;
    wire [31:0] _5027;
    wire [31:0] _5028;
    wire [31:0] _5029;
    wire _5030;
    wire [31:0] _5031;
    wire _5032;
    wire [31:0] _5033;
    wire [31:0] _2658;
    reg [31:0] _2660;
    wire [31:0] _3289;
    wire _3294;
    wire _3295;
    wire _3296;
    wire [31:0] _3316;
    wire _3298;
    wire _3299;
    wire _3300;
    wire _3311;
    wire _3319;
    wire _3313;
    wire _3315;
    wire _3321;
    wire _3323;
    wire [31:0] _3324;
    wire [31:0] _3379;
    reg [31:0] _3381;
    wire [31:0] _3384 = 32'b00000000000000000000000000000000;
    wire [31:0] _3382 = 32'b00000000000000000000000000000000;
    wire _4569;
    wire _4570;
    wire _4571;
    wire _4572;
    wire _4573;
    wire _4574;
    wire _4575;
    wire _4576;
    wire _4577;
    wire _4578;
    wire _4579;
    wire _4580;
    wire _4581;
    wire _4582;
    wire _4583;
    wire _4584;
    wire _4585;
    wire _4586;
    wire _4587;
    wire _4588;
    wire _4589;
    wire _4590;
    wire _4591;
    wire _4592;
    wire _4593;
    wire _4594;
    wire _4595;
    wire _4596;
    wire _4597;
    wire _4598;
    wire _4599;
    wire _4600;
    wire _4601;
    wire _4602;
    wire _4603;
    wire _4604;
    wire _4605;
    wire _4606;
    wire _4607;
    wire _4608;
    wire _4609;
    wire _4610;
    wire _4611;
    wire _4612;
    wire _4613;
    wire _4614;
    wire _4615;
    wire _4616;
    wire _4617;
    wire _4618;
    wire _4619;
    wire _4620;
    wire _4621;
    wire _4622;
    wire _4623;
    wire _4624;
    wire _4625;
    wire _4626;
    wire _4627;
    wire _4628;
    wire _4629;
    wire _4630;
    wire _4631;
    wire [31:0] _4632;
    wire [31:0] _4633;
    wire [31:0] _4634;
    wire [31:0] _4635;
    wire [31:0] _4636;
    wire [31:0] _4637;
    wire [31:0] _3767;
    wire [63:0] _3344 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3342 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3961 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _3962;
    wire [63:0] _4872;
    wire [63:0] _3343;
    reg [63:0] count_cycle;
    wire [31:0] _3765;
    wire [31:0] _3771;
    wire [31:0] _3763;
    wire [63:0] _3340 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3338 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3549 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _3550;
    wire [63:0] _4873;
    wire [63:0] _4874;
    wire [63:0] _4875;
    wire [63:0] _4876;
    wire _4877;
    wire [63:0] _4878;
    wire [63:0] _3339;
    reg [63:0] _3341;
    wire [31:0] _3761;
    wire _3764;
    wire [31:0] _3769;
    wire _3766;
    wire _3768;
    wire _3772;
    wire [31:0] _3773;
    wire [31:0] _4638;
    wire [31:0] _4639;
    wire [31:0] _4640;
    wire [31:0] _4641;
    wire [31:0] _4642;
    wire [31:0] _4643;
    wire [31:0] _4644;
    wire [31:0] _4645;
    wire [31:0] _4646;
    wire [31:0] _4647;
    wire [31:0] _3374 = 32'b00000000000000000000000000000000;
    wire [31:0] _39 = 32'b00000000000000000000000000000000;
    wire _4668;
    wire [31:0] _4669;
    wire [31:0] _3373;
    reg [31:0] _3375;
    wire [31:0] _3814;
    wire [31:0] _4648;
    wire [15:0] _3902;
    wire _3903;
    wire [1:0] _3904;
    wire [3:0] _3905;
    wire [7:0] _3906;
    wire [15:0] _3907;
    wire [31:0] _3909;
    wire [31:0] _3910;
    wire [7:0] _3893;
    wire _3894;
    wire [1:0] _3895;
    wire [3:0] _3896;
    wire [7:0] _3897;
    wire [15:0] _3898;
    wire [23:0] _3899;
    wire [31:0] _3901;
    wire _3364 = 1'b0;
    wire _3362 = 1'b0;
    wire _3656 = 1'b0;
    wire _3919;
    wire _4746;
    wire _4747;
    wire _4748;
    wire _4749;
    wire _4750;
    wire _4751;
    wire _3363;
    reg _3365;
    wire _3368 = 1'b0;
    wire _3366 = 1'b0;
    wire _3657 = 1'b0;
    wire _3920;
    wire _4740;
    wire _4741;
    wire _4742;
    wire _4743;
    wire _4744;
    wire _4745;
    wire _3367;
    reg _3369;
    wire _3911;
    wire [31:0] _3912;
    wire _3914;
    wire _3915;
    wire [31:0] _4649;
    wire [31:0] _4650;
    wire [31:0] _4130 = 32'b00000000000000000000000000000000;
    wire _4651;
    wire [31:0] _4652;
    wire _4653;
    wire [31:0] _4654;
    wire _4655;
    wire [31:0] _4656;
    wire _4657;
    wire [31:0] _4658;
    wire _4659;
    wire [31:0] _4660;
    wire _4661;
    wire [31:0] _4662;
    wire [31:0] _3383;
    reg [31:0] _3385;
    wire _3352 = 1'b0;
    wire _3350 = 1'b0;
    wire _3659 = 1'b0;
    wire _3807 = 1'b1;
    wire _4850;
    wire _4851;
    wire _4852;
    wire _4853;
    wire _4854;
    wire _3351;
    reg _3353;
    wire [31:0] _3675;
    wire [31:0] _3676;
    wire [31:0] _40 = 32'b00000000000000000000000000010000;
    wire [31:0] _4663;
    wire [31:0] _4664;
    wire [31:0] _4665;
    wire [31:0] _3376 = 32'b00000000000000000000000000000000;
    wire _4666;
    wire [31:0] _4667;
    wire [31:0] _3377;
    wire [31:0] _4735;
    wire [31:0] _4736;
    wire [31:0] _4737;
    wire _4738;
    wire [31:0] _4739;
    wire [31:0] _3370;
    reg [31:0] _3372;
    wire [31:0] _4970;
    wire [31:0] _3662;
    wire [31:0] _3663;
    wire [31:0] _4971;
    wire [31:0] _4972;
    wire [31:0] _4973;
    wire [31:0] _4974;
    wire _3348 = 1'b0;
    wire _3346 = 1'b0;
    wire _3545 = 1'b1;
    wire _3548;
    wire _4855;
    wire _3658 = 1'b0;
    wire _4856;
    wire _3558;
    wire _3336 = 1'b0;
    wire _3334 = 1'b0;
    wire _3553 = 1'b1;
    wire _4879;
    wire _4880;
    wire _4881;
    wire _4882;
    wire _4883;
    wire _4884;
    wire _4885;
    wire _4886;
    wire _4887;
    wire _4888;
    wire _4889;
    wire _4890;
    wire _4891;
    wire _4892;
    wire _4893;
    wire _4894;
    wire _4895;
    wire _4896;
    wire _4897;
    wire _4898;
    wire _4899;
    wire _4900;
    wire _4901;
    wire _4902;
    wire _4903;
    wire _4904;
    wire _4905;
    wire _4906;
    wire _4907;
    wire _4908;
    wire _4909;
    wire [31:0] _3400 = 32'b00000000000000000000000000000000;
    wire [31:0] _3398 = 32'b00000000000000000000000000000000;
    wire _3436 = 1'b0;
    wire _3705;
    wire _4466;
    wire _4467;
    wire _4468;
    wire _4469;
    wire _4470;
    wire _4471;
    wire _4472;
    wire _4473;
    wire _4474;
    wire _4475;
    wire _3435;
    reg _3437;
    wire _3442 = 1'b0;
    wire _3707;
    wire _4446;
    wire _4447;
    wire _4448;
    wire _4449;
    wire _4450;
    wire _4451;
    wire _4452;
    wire _4453;
    wire _4454;
    wire _4455;
    wire _3441;
    reg _3443;
    wire _3445 = 1'b0;
    wire _3708;
    wire _4436;
    wire _4437;
    wire _4438;
    wire _4439;
    wire _4440;
    wire _4441;
    wire _4442;
    wire _4443;
    wire _4444;
    wire _4445;
    wire _3444;
    reg _3446;
    wire _3448 = 1'b0;
    wire _3709;
    wire _4426;
    wire _4427;
    wire _4428;
    wire _4429;
    wire _4430;
    wire _4431;
    wire _4432;
    wire _4433;
    wire _4434;
    wire _4435;
    wire _3447;
    reg _3449;
    wire _3451 = 1'b0;
    wire _3710;
    wire _4416;
    wire _4417;
    wire _4418;
    wire _4419;
    wire _4420;
    wire _4421;
    wire _4422;
    wire _4423;
    wire _4424;
    wire _4425;
    wire _3450;
    reg _3452;
    wire _3454 = 1'b0;
    wire _3711;
    wire _4406;
    wire _4407;
    wire _4408;
    wire _4409;
    wire _4410;
    wire _4411;
    wire _4412;
    wire _4413;
    wire _4414;
    wire _4415;
    wire _3453;
    reg _3455;
    wire _3457 = 1'b0;
    wire _3712;
    wire _4396;
    wire _4397;
    wire _4398;
    wire _4399;
    wire _4400;
    wire _4401;
    wire _4402;
    wire _4403;
    wire _4404;
    wire _4405;
    wire _3456;
    reg _3458;
    wire _3460 = 1'b0;
    wire _3713;
    wire _4386;
    wire _4387;
    wire _4388;
    wire _4389;
    wire _4390;
    wire _4391;
    wire _4392;
    wire _4393;
    wire _4394;
    wire _4395;
    wire _3459;
    reg _3461;
    wire _3463 = 1'b0;
    wire _3714;
    wire _4376;
    wire _4377;
    wire _4378;
    wire _4379;
    wire _4380;
    wire _4381;
    wire _4382;
    wire _4383;
    wire _4384;
    wire _4385;
    wire _3462;
    reg _3464;
    wire _3466 = 1'b0;
    wire _3715;
    wire _4366;
    wire _4367;
    wire _4368;
    wire _4369;
    wire _4370;
    wire _4371;
    wire _4372;
    wire _4373;
    wire _4374;
    wire _4375;
    wire _3465;
    reg _3467;
    wire _3469 = 1'b0;
    wire _3716;
    wire _4356;
    wire _4357;
    wire _4358;
    wire _4359;
    wire _4360;
    wire _4361;
    wire _4362;
    wire _4363;
    wire _4364;
    wire _4365;
    wire _3468;
    reg _3470;
    wire _3472 = 1'b0;
    wire _3717;
    wire _4346;
    wire _4347;
    wire _4348;
    wire _4349;
    wire _4350;
    wire _4351;
    wire _4352;
    wire _4353;
    wire _4354;
    wire _4355;
    wire _3471;
    reg _3473;
    wire _3475 = 1'b0;
    wire _3718;
    wire _4336;
    wire _4337;
    wire _4338;
    wire _4339;
    wire _4340;
    wire _4341;
    wire _4342;
    wire _4343;
    wire _4344;
    wire _4345;
    wire _3474;
    reg _3476;
    wire _3478 = 1'b0;
    wire _3719;
    wire _4326;
    wire _4327;
    wire _4328;
    wire _4329;
    wire _4330;
    wire _4331;
    wire _4332;
    wire _4333;
    wire _4334;
    wire _4335;
    wire _3477;
    reg _3479;
    wire _3481 = 1'b0;
    wire _3720;
    wire _4316;
    wire _4317;
    wire _4318;
    wire _4319;
    wire _4320;
    wire _4321;
    wire _4322;
    wire _4323;
    wire _4324;
    wire _4325;
    wire _3480;
    reg _3482;
    wire _3484 = 1'b0;
    wire _3721;
    wire _4306;
    wire _4307;
    wire _4308;
    wire _4309;
    wire _4310;
    wire _4311;
    wire _4312;
    wire _4313;
    wire _4314;
    wire _4315;
    wire _3483;
    reg _3485;
    wire _3487 = 1'b0;
    wire _3722;
    wire _4296;
    wire _4297;
    wire _4298;
    wire _4299;
    wire _4300;
    wire _4301;
    wire _4302;
    wire _4303;
    wire _4304;
    wire _4305;
    wire _3486;
    reg _3488;
    wire _3490 = 1'b0;
    wire _3723;
    wire _4286;
    wire _4287;
    wire _4288;
    wire _4289;
    wire _4290;
    wire _4291;
    wire _4292;
    wire _4293;
    wire _4294;
    wire _4295;
    wire _3489;
    reg _3491;
    wire _3493 = 1'b0;
    wire _3724;
    wire _4276;
    wire _4277;
    wire _4278;
    wire _4279;
    wire _4280;
    wire _4281;
    wire _4282;
    wire _4283;
    wire _4284;
    wire _4285;
    wire _3492;
    reg _3494;
    wire _3496 = 1'b0;
    wire _3725;
    wire _4266;
    wire _4267;
    wire _4268;
    wire _4269;
    wire _4270;
    wire _4271;
    wire _4272;
    wire _4273;
    wire _4274;
    wire _4275;
    wire _3495;
    reg _3497;
    wire _3499 = 1'b0;
    wire _3726;
    wire _4256;
    wire _4257;
    wire _4258;
    wire _4259;
    wire _4260;
    wire _4261;
    wire _4262;
    wire _4263;
    wire _4264;
    wire _4265;
    wire _3498;
    reg _3500;
    wire _3502 = 1'b0;
    wire _3727;
    wire _4246;
    wire _4247;
    wire _4248;
    wire _4249;
    wire _4250;
    wire _4251;
    wire _4252;
    wire _4253;
    wire _4254;
    wire _4255;
    wire _3501;
    reg _3503;
    wire _3505 = 1'b0;
    wire _3728;
    wire _4236;
    wire _4237;
    wire _4238;
    wire _4239;
    wire _4240;
    wire _4241;
    wire _4242;
    wire _4243;
    wire _4244;
    wire _4245;
    wire _3504;
    reg _3506;
    wire _3508 = 1'b0;
    wire _3729;
    wire _4226;
    wire _4227;
    wire _4228;
    wire _4229;
    wire _4230;
    wire _4231;
    wire _4232;
    wire _4233;
    wire _4234;
    wire _4235;
    wire _3507;
    reg _3509;
    wire _3511 = 1'b0;
    wire _3730;
    wire _4216;
    wire _4217;
    wire _4218;
    wire _4219;
    wire _4220;
    wire _4221;
    wire _4222;
    wire _4223;
    wire _4224;
    wire _4225;
    wire _3510;
    reg _3512;
    wire _3514 = 1'b0;
    wire _3731;
    wire _4206;
    wire _4207;
    wire _4208;
    wire _4209;
    wire _4210;
    wire _4211;
    wire _4212;
    wire _4213;
    wire _4214;
    wire _4215;
    wire _3513;
    reg _3515;
    wire _3517 = 1'b0;
    wire _3732;
    wire _4196;
    wire _4197;
    wire _4198;
    wire _4199;
    wire _4200;
    wire _4201;
    wire _4202;
    wire _4203;
    wire _4204;
    wire _4205;
    wire _3516;
    reg _3518;
    wire _3520 = 1'b0;
    wire _3733;
    wire _4186;
    wire _4187;
    wire _4188;
    wire _4189;
    wire _4190;
    wire _4191;
    wire _4192;
    wire _4193;
    wire _4194;
    wire _4195;
    wire _3519;
    reg _3521;
    wire _3523 = 1'b0;
    wire _3734;
    wire _4176;
    wire _4177;
    wire _4178;
    wire _4179;
    wire _4180;
    wire _4181;
    wire _4182;
    wire _4183;
    wire _4184;
    wire _4185;
    wire _3522;
    reg _3524;
    wire _3526 = 1'b0;
    wire _3735;
    wire _4166;
    wire _4167;
    wire _4168;
    wire _4169;
    wire _4170;
    wire _4171;
    wire _4172;
    wire _4173;
    wire _4174;
    wire _4175;
    wire _3525;
    reg _3527;
    wire _3529 = 1'b0;
    wire _3736;
    wire _4156;
    wire _4157;
    wire _4158;
    wire _4159;
    wire _4160;
    wire _4161;
    wire _4162;
    wire _4163;
    wire _4164;
    wire _4165;
    wire _3528;
    reg _3530;
    wire [31:0] _3531;
    wire [31:0] _3661;
    wire [31:0] _4525;
    wire [31:0] _4526;
    wire [31:0] _4527;
    wire [31:0] _4528;
    wire _3951 = 1'b1;
    wire [31:0] _3954 = 32'b00000000000000000000000000000000;
    wire [31:0] _3952 = 32'b00000000000000000000000000000001;
    wire [31:0] _3953;
    wire _3955;
    wire _4523;
    wire _3970;
    wire _3971;
    wire _3972;
    wire _3973;
    wire _3974;
    wire _4522;
    wire [31:0] _3956 = 32'b00000000000000000000000000000000;
    wire [31:0] _3537 = 32'b00000000000000000000000000000000;
    wire [31:0] _3535 = 32'b00000000000000000000000000000000;
    wire _3701;
    wire _3702;
    wire _3703;
    wire [31:0] _4134;
    wire [31:0] _4135;
    wire [31:0] _4136;
    wire [31:0] _4137;
    wire [31:0] _4138;
    wire [31:0] _4139;
    wire [31:0] _4140;
    wire [31:0] _4141;
    wire [31:0] _3949 = 32'b00000000000000000000000000000001;
    wire [31:0] _3950;
    wire [31:0] _4133;
    wire _4142;
    wire [31:0] _4143;
    wire [31:0] _3536;
    reg [31:0] _3538;
    wire _3957;
    wire _3958;
    wire _3959;
    wire _3960;
    wire _4524;
    wire _3402;
    wire _3781 = 1'b1;
    wire _3782;
    wire _3783;
    wire _3784;
    wire _3785;
    wire _4507;
    wire _4508;
    wire _4509;
    wire _4510;
    wire _3776 = 1'b1;
    wire _3777;
    wire _3778;
    wire _3779;
    wire _3780;
    wire _4511;
    wire _4512;
    wire _4513;
    wire _3796 = 1'b1;
    wire _3396 = 1'b0;
    wire _3394 = 1'b0;
    wire _3669 = 1'b1;
    wire _4531;
    wire _4532;
    wire _4533;
    wire _3742 = 1'b0;
    wire _4534;
    wire _4535;
    wire _4536;
    wire _4537;
    wire _4538;
    wire _4539;
    wire _4540;
    wire _4541;
    wire _4542;
    wire _4543;
    wire _3395;
    reg _3397;
    wire _3797;
    wire _3439 = 1'b0;
    wire [31:0] _37 = 32'b00000000000000000000000000000000;
    wire _3241;
    wire _3242;
    wire [31:0] _3244 = 32'b00000000000000000000000000000000;
    wire [31:0] _3243 = 32'b00000000000000000000000000000000;
    reg [31:0] _3245;
    wire _3236;
    wire _3237;
    wire [31:0] _3239 = 32'b00000000000000000000000000000000;
    wire [31:0] _3238 = 32'b00000000000000000000000000000000;
    reg [31:0] _3240;
    wire _3231;
    wire _3232;
    wire [31:0] _3234 = 32'b00000000000000000000000000000000;
    wire [31:0] _3233 = 32'b00000000000000000000000000000000;
    reg [31:0] _3235;
    wire _3226;
    wire _3227;
    wire [31:0] _3229 = 32'b00000000000000000000000000000000;
    wire [31:0] _3228 = 32'b00000000000000000000000000000000;
    reg [31:0] _3230;
    wire _3221;
    wire _3222;
    wire [31:0] _3224 = 32'b00000000000000000000000000000000;
    wire [31:0] _3223 = 32'b00000000000000000000000000000000;
    reg [31:0] _3225;
    wire _3216;
    wire _3217;
    wire [31:0] _3219 = 32'b00000000000000000000000000000000;
    wire [31:0] _3218 = 32'b00000000000000000000000000000000;
    reg [31:0] _3220;
    wire _3211;
    wire _3212;
    wire [31:0] _3214 = 32'b00000000000000000000000000000000;
    wire [31:0] _3213 = 32'b00000000000000000000000000000000;
    reg [31:0] _3215;
    wire _3206;
    wire _3207;
    wire [31:0] _3209 = 32'b00000000000000000000000000000000;
    wire [31:0] _3208 = 32'b00000000000000000000000000000000;
    reg [31:0] _3210;
    wire _3201;
    wire _3202;
    wire [31:0] _3204 = 32'b00000000000000000000000000000000;
    wire [31:0] _3203 = 32'b00000000000000000000000000000000;
    reg [31:0] _3205;
    wire _3196;
    wire _3197;
    wire [31:0] _3199 = 32'b00000000000000000000000000000000;
    wire [31:0] _3198 = 32'b00000000000000000000000000000000;
    reg [31:0] _3200;
    wire _3191;
    wire _3192;
    wire [31:0] _3194 = 32'b00000000000000000000000000000000;
    wire [31:0] _3193 = 32'b00000000000000000000000000000000;
    reg [31:0] _3195;
    wire _3186;
    wire _3187;
    wire [31:0] _3189 = 32'b00000000000000000000000000000000;
    wire [31:0] _3188 = 32'b00000000000000000000000000000000;
    reg [31:0] _3190;
    wire _3181;
    wire _3182;
    wire [31:0] _3184 = 32'b00000000000000000000000000000000;
    wire [31:0] _3183 = 32'b00000000000000000000000000000000;
    reg [31:0] _3185;
    wire _3176;
    wire _3177;
    wire [31:0] _3179 = 32'b00000000000000000000000000000000;
    wire [31:0] _3178 = 32'b00000000000000000000000000000000;
    reg [31:0] _3180;
    wire _3171;
    wire _3172;
    wire [31:0] _3174 = 32'b00000000000000000000000000000000;
    wire [31:0] _3173 = 32'b00000000000000000000000000000000;
    reg [31:0] _3175;
    wire _3166;
    wire _3167;
    wire [31:0] _3169 = 32'b00000000000000000000000000000000;
    wire [31:0] _3168 = 32'b00000000000000000000000000000000;
    reg [31:0] _3170;
    wire _3161;
    wire _3162;
    wire [31:0] _3164 = 32'b00000000000000000000000000000000;
    wire [31:0] _3163 = 32'b00000000000000000000000000000000;
    reg [31:0] _3165;
    wire _3156;
    wire _3157;
    wire [31:0] _3159 = 32'b00000000000000000000000000000000;
    wire [31:0] _3158 = 32'b00000000000000000000000000000000;
    reg [31:0] _3160;
    wire _3151;
    wire _3152;
    wire [31:0] _3154 = 32'b00000000000000000000000000000000;
    wire [31:0] _3153 = 32'b00000000000000000000000000000000;
    reg [31:0] _3155;
    wire _3146;
    wire _3147;
    wire [31:0] _3149 = 32'b00000000000000000000000000000000;
    wire [31:0] _3148 = 32'b00000000000000000000000000000000;
    reg [31:0] _3150;
    wire _3141;
    wire _3142;
    wire [31:0] _3144 = 32'b00000000000000000000000000000000;
    wire [31:0] _3143 = 32'b00000000000000000000000000000000;
    reg [31:0] _3145;
    wire _3136;
    wire _3137;
    wire [31:0] _3139 = 32'b00000000000000000000000000000000;
    wire [31:0] _3138 = 32'b00000000000000000000000000000000;
    reg [31:0] _3140;
    wire _3131;
    wire _3132;
    wire [31:0] _3134 = 32'b00000000000000000000000000000000;
    wire [31:0] _3133 = 32'b00000000000000000000000000000000;
    reg [31:0] _3135;
    wire _3126;
    wire _3127;
    wire [31:0] _3129 = 32'b00000000000000000000000000000000;
    wire [31:0] _3128 = 32'b00000000000000000000000000000000;
    reg [31:0] _3130;
    wire _3121;
    wire _3122;
    wire [31:0] _3124 = 32'b00000000000000000000000000000000;
    wire [31:0] _3123 = 32'b00000000000000000000000000000000;
    reg [31:0] _3125;
    wire _3116;
    wire _3117;
    wire [31:0] _3119 = 32'b00000000000000000000000000000000;
    wire [31:0] _3118 = 32'b00000000000000000000000000000000;
    reg [31:0] _3120;
    wire _3111;
    wire _3112;
    wire [31:0] _3114 = 32'b00000000000000000000000000000000;
    wire [31:0] _3113 = 32'b00000000000000000000000000000000;
    reg [31:0] _3115;
    wire _3106;
    wire _3107;
    wire [31:0] _3109 = 32'b00000000000000000000000000000000;
    wire [31:0] _3108 = 32'b00000000000000000000000000000000;
    reg [31:0] _3110;
    wire _3101;
    wire _3102;
    wire [31:0] _3104 = 32'b00000000000000000000000000000000;
    wire [31:0] _3103 = 32'b00000000000000000000000000000000;
    reg [31:0] _3105;
    wire _3096;
    wire _3097;
    wire [31:0] _3099 = 32'b00000000000000000000000000000000;
    wire [31:0] _3098 = 32'b00000000000000000000000000000000;
    reg [31:0] _3100;
    wire _3091;
    wire _3092;
    wire [31:0] _3094 = 32'b00000000000000000000000000000000;
    wire [31:0] _3093 = 32'b00000000000000000000000000000000;
    reg [31:0] _3095;
    wire _3086;
    wire _3087;
    wire [31:0] _3089 = 32'b00000000000000000000000000000000;
    wire [31:0] _3088 = 32'b00000000000000000000000000000000;
    reg [31:0] _3090;
    wire _3081;
    wire _3082;
    wire [31:0] _3084 = 32'b00000000000000000000000000000000;
    wire [31:0] _3083 = 32'b00000000000000000000000000000000;
    reg [31:0] _3085;
    wire _3076;
    wire _3077;
    wire [31:0] _3079 = 32'b00000000000000000000000000000000;
    wire [31:0] _3078 = 32'b00000000000000000000000000000000;
    reg [31:0] _3080;
    wire _2682;
    wire _2685;
    wire _2693;
    wire _2713;
    wire _2761;
    wire _2873;
    wire _2683;
    wire _2684;
    wire _2692;
    wire _2712;
    wire _2760;
    wire _2872;
    wire _2686;
    wire _2688;
    wire _2691;
    wire _2711;
    wire _2759;
    wire _2871;
    wire _2687;
    wire _2689;
    wire _2690;
    wire _2710;
    wire _2758;
    wire _2870;
    wire _2694;
    wire _2697;
    wire _2704;
    wire _2709;
    wire _2757;
    wire _2869;
    wire _2695;
    wire _2696;
    wire _2703;
    wire _2708;
    wire _2756;
    wire _2868;
    wire _2698;
    wire _2700;
    wire _2702;
    wire _2707;
    wire _2755;
    wire _2867;
    wire _2699;
    wire _2701;
    wire _2705;
    wire _2706;
    wire _2754;
    wire _2866;
    wire _2714;
    wire _2717;
    wire _2725;
    wire _2744;
    wire _2753;
    wire _2865;
    wire _2715;
    wire _2716;
    wire _2724;
    wire _2743;
    wire _2752;
    wire _2864;
    wire _2718;
    wire _2720;
    wire _2723;
    wire _2742;
    wire _2751;
    wire _2863;
    wire _2719;
    wire _2721;
    wire _2722;
    wire _2741;
    wire _2750;
    wire _2862;
    wire _2726;
    wire _2729;
    wire _2736;
    wire _2740;
    wire _2749;
    wire _2861;
    wire _2727;
    wire _2728;
    wire _2735;
    wire _2739;
    wire _2748;
    wire _2860;
    wire _2730;
    wire _2732;
    wire _2734;
    wire _2738;
    wire _2747;
    wire _2859;
    wire _2731;
    wire _2733;
    wire _2737;
    wire _2745;
    wire _2746;
    wire _2858;
    wire _2762;
    wire _2765;
    wire _2773;
    wire _2793;
    wire _2840;
    wire _2857;
    wire _2763;
    wire _2764;
    wire _2772;
    wire _2792;
    wire _2839;
    wire _2856;
    wire _2766;
    wire _2768;
    wire _2771;
    wire _2791;
    wire _2838;
    wire _2855;
    wire _2767;
    wire _2769;
    wire _2770;
    wire _2790;
    wire _2837;
    wire _2854;
    wire _2774;
    wire _2777;
    wire _2784;
    wire _2789;
    wire _2836;
    wire _2853;
    wire _2775;
    wire _2776;
    wire _2783;
    wire _2788;
    wire _2835;
    wire _2852;
    wire _2778;
    wire _2780;
    wire _2782;
    wire _2787;
    wire _2834;
    wire _2851;
    wire _2779;
    wire _2781;
    wire _2785;
    wire _2786;
    wire _2833;
    wire _2850;
    wire _2794;
    wire _2797;
    wire _2805;
    wire _2824;
    wire _2832;
    wire _2849;
    wire _2795;
    wire _2796;
    wire _2804;
    wire _2823;
    wire _2831;
    wire _2848;
    wire _2798;
    wire _2800;
    wire _2803;
    wire _2822;
    wire _2830;
    wire _2847;
    wire _2799;
    wire _2801;
    wire _2802;
    wire _2821;
    wire _2829;
    wire _2846;
    wire _2806;
    wire _2809;
    wire _2816;
    wire _2820;
    wire _2828;
    wire _2845;
    wire _2807;
    wire _2808;
    wire _2815;
    wire _2819;
    wire _2827;
    wire _2844;
    wire _2810;
    wire _2812;
    wire _2814;
    wire _2818;
    wire _2826;
    wire _2843;
    wire _2811;
    wire _2813;
    wire _2817;
    wire _2825;
    wire _2841;
    wire _2842;
    wire _2874;
    wire _2877;
    wire _2885;
    wire _2905;
    wire _2953;
    wire _3064;
    wire _2875;
    wire _2876;
    wire _2884;
    wire _2904;
    wire _2952;
    wire _3063;
    wire _2878;
    wire _2880;
    wire _2883;
    wire _2903;
    wire _2951;
    wire _3062;
    wire _2879;
    wire _2881;
    wire _2882;
    wire _2902;
    wire _2950;
    wire _3061;
    wire _2886;
    wire _2889;
    wire _2896;
    wire _2901;
    wire _2949;
    wire _3060;
    wire _2887;
    wire _2888;
    wire _2895;
    wire _2900;
    wire _2948;
    wire _3059;
    wire _2890;
    wire _2892;
    wire _2894;
    wire _2899;
    wire _2947;
    wire _3058;
    wire _2891;
    wire _2893;
    wire _2897;
    wire _2898;
    wire _2946;
    wire _3057;
    wire _2906;
    wire _2909;
    wire _2917;
    wire _2936;
    wire _2945;
    wire _3056;
    wire _2907;
    wire _2908;
    wire _2916;
    wire _2935;
    wire _2944;
    wire _3055;
    wire _2910;
    wire _2912;
    wire _2915;
    wire _2934;
    wire _2943;
    wire _3054;
    wire _2911;
    wire _2913;
    wire _2914;
    wire _2933;
    wire _2942;
    wire _3053;
    wire _2918;
    wire _2921;
    wire _2928;
    wire _2932;
    wire _2941;
    wire _3052;
    wire _2919;
    wire _2920;
    wire _2927;
    wire _2931;
    wire _2940;
    wire _3051;
    wire _2922;
    wire _2924;
    wire _2926;
    wire _2930;
    wire _2939;
    wire _3050;
    wire _2923;
    wire _2925;
    wire _2929;
    wire _2937;
    wire _2938;
    wire _3049;
    wire _2954;
    wire _2957;
    wire _2965;
    wire _2985;
    wire _3032;
    wire _3048;
    wire _2955;
    wire _2956;
    wire _2964;
    wire _2984;
    wire _3031;
    wire _3047;
    wire _2958;
    wire _2960;
    wire _2963;
    wire _2983;
    wire _3030;
    wire _3046;
    wire _2959;
    wire _2961;
    wire _2962;
    wire _2982;
    wire _3029;
    wire _3045;
    wire _2966;
    wire _2969;
    wire _2976;
    wire _2981;
    wire _3028;
    wire _3044;
    wire _2967;
    wire _2968;
    wire _2975;
    wire _2980;
    wire _3027;
    wire _3043;
    wire _2970;
    wire _2972;
    wire _2974;
    wire _2979;
    wire _3026;
    wire _3042;
    wire _2971;
    wire _2973;
    wire _2977;
    wire _2978;
    wire _3025;
    wire _3041;
    wire _2986;
    wire _2989;
    wire _2997;
    wire _3016;
    wire _3024;
    wire _3040;
    wire _2987;
    wire _2988;
    wire _2996;
    wire _3015;
    wire _3023;
    wire _3039;
    wire _2990;
    wire _2992;
    wire _2995;
    wire _3014;
    wire _3022;
    wire _3038;
    wire _2991;
    wire _2993;
    wire _2994;
    wire _3013;
    wire _3021;
    wire _3037;
    wire _2998;
    wire _3001;
    wire _3008;
    wire _3012;
    wire _3020;
    wire _3036;
    wire _2999;
    wire _3000;
    wire _3007;
    wire _3011;
    wire _3019;
    wire _3035;
    wire _3002;
    wire _3004;
    wire _3006;
    wire _3010;
    wire _3018;
    wire _3034;
    wire _2676;
    wire _2677;
    wire _3003;
    wire _2678;
    wire _3005;
    wire _2679;
    wire _3009;
    wire _2680;
    wire _3017;
    wire [5:0] _2671 = 6'b000000;
    wire [5:0] _2669 = 6'b000000;
    wire _3565;
    wire [4:0] _3568 = 5'b00000;
    wire [5:0] _3570;
    wire [5:0] _3571 = 6'b100000;
    wire [5:0] _3572;
    wire [5:0] _3563 = 6'b000100;
    wire [5:0] _3562 = 6'b000011;
    wire _3564;
    wire [5:0] _4978;
    wire [5:0] _4979;
    wire [5:0] _4980;
    wire [5:0] _3747 = 6'b100000;
    wire [5:0] _3748;
    wire [5:0] _4981;
    wire [5:0] _4982;
    wire [5:0] _4983;
    wire [5:0] _4984;
    wire [5:0] _4985;
    wire [5:0] _3812 = 6'b000000;
    wire [5:0] _4986;
    wire _4987;
    wire [5:0] _4988;
    wire _4989;
    wire [5:0] _4990;
    wire _4991;
    wire [5:0] _4992;
    wire [5:0] _2670;
    reg [5:0] _2672;
    wire _2681;
    wire _3033;
    wire [63:0] _3065;
    wire _3071;
    wire _4958;
    wire _4959;
    wire _4960;
    wire _4961;
    wire _3666;
    wire _3667;
    wire _4962;
    wire [1:0] _3392 = 2'b00;
    wire [1:0] _3390 = 2'b00;
    wire [1:0] _3578 = 2'b01;
    wire [1:0] _3574 = 2'b10;
    wire [1:0] _3573 = 2'b00;
    wire [1:0] _3575 = 2'b01;
    wire _3576;
    wire [1:0] _3577;
    wire [1:0] _3579 = 2'b00;
    wire _3580;
    wire [1:0] _3581;
    wire [1:0] _4544;
    wire _4545;
    wire [1:0] _4546;
    wire [1:0] _3391;
    reg [1:0] _3393;
    wire _3670;
    wire _3671;
    wire _4963;
    wire _4964;
    wire _4965;
    wire _4966;
    wire _4967;
    wire _2675;
    wire _3072;
    wire [31:0] _3074 = 32'b00000000000000000000000000000000;
    wire [31:0] _3073 = 32'b00000000000000000000000000000000;
    reg [31:0] _3075;
    reg [31:0] _3247;
    wire [31:0] _3681 = 32'b00000000000000000000000000000000;
    wire [5:0] _3682 = 6'b000000;
    wire _3683;
    wire _3684;
    wire [31:0] _3685;
    wire [31:0] _3704;
    wire _3706;
    wire _4456;
    wire _3738;
    wire _3739;
    wire _4457;
    wire _4458;
    wire _4459;
    wire _4460;
    wire _4461;
    wire _4462;
    wire _4463;
    wire _4464;
    wire _4465;
    wire _3438;
    reg _3440;
    wire _3798;
    wire _3799;
    wire _3800;
    wire _4514;
    wire _3328 = 1'b0;
    wire _3326 = 1'b0;
    wire [3:0] _3963 = 4'b0000;
    wire [3:0] _3332 = 4'b0000;
    wire [3:0] _3330 = 4'b0000;
    wire [3:0] _3966 = 4'b0001;
    wire [3:0] _3967;
    wire _4947;
    wire _4948;
    wire _4949;
    wire _4950;
    wire _4951;
    wire _4952;
    wire _4953;
    wire [3:0] _4954;
    wire [3:0] _3965 = 4'b1111;
    wire _3968;
    wire _2631 = 1'b0;
    wire _2629 = 1'b0;
    wire _3786 = 1'b0;
    wire _3789 = 1'b1;
    wire _5160;
    wire _5161;
    wire _5162;
    wire _5163;
    wire _3801 = 1'b0;
    wire _3803 = 1'b1;
    wire _5164;
    wire _5165;
    wire _5166;
    wire _5167;
    wire _5168;
    wire _5169;
    wire _2630;
    reg _2632;
    wire _3969;
    wire [3:0] _4955;
    wire [3:0] _4956;
    wire [3:0] _3331;
    reg [3:0] _3333;
    wire _3964;
    wire _4957;
    wire _3327;
    reg _3329;
    wire _4515;
    wire _4516;
    wire _3804;
    wire _3805;
    wire _4517;
    wire _3975;
    wire _3976;
    wire _3977;
    wire _3978;
    wire _3979;
    wire _4506;
    wire _4518;
    wire _4519;
    wire _4520;
    wire _4521;
    wire _3403;
    wire _3980;
    wire _3981;
    wire _3982;
    wire _3983;
    wire _3984;
    wire _4505;
    wire _3404;
    wire _3985;
    wire _3986;
    wire _3987;
    wire _3988;
    wire _3989;
    wire _4504;
    wire _3405;
    wire _3990;
    wire _3991;
    wire _3992;
    wire _3993;
    wire _3994;
    wire _4503;
    wire _3406;
    wire _3995;
    wire _3996;
    wire _3997;
    wire _3998;
    wire _3999;
    wire _4502;
    wire _3407;
    wire _4000;
    wire _4001;
    wire _4002;
    wire _4003;
    wire _4004;
    wire _4501;
    wire _3408;
    wire _4005;
    wire _4006;
    wire _4007;
    wire _4008;
    wire _4009;
    wire _4500;
    wire _3409;
    wire _4010;
    wire _4011;
    wire _4012;
    wire _4013;
    wire _4014;
    wire _4499;
    wire _3410;
    wire _4015;
    wire _4016;
    wire _4017;
    wire _4018;
    wire _4019;
    wire _4498;
    wire _3411;
    wire _4020;
    wire _4021;
    wire _4022;
    wire _4023;
    wire _4024;
    wire _4497;
    wire _3412;
    wire _4025;
    wire _4026;
    wire _4027;
    wire _4028;
    wire _4029;
    wire _4496;
    wire _3413;
    wire _4030;
    wire _4031;
    wire _4032;
    wire _4033;
    wire _4034;
    wire _4495;
    wire _3414;
    wire _4035;
    wire _4036;
    wire _4037;
    wire _4038;
    wire _4039;
    wire _4494;
    wire _3415;
    wire _4040;
    wire _4041;
    wire _4042;
    wire _4043;
    wire _4044;
    wire _4493;
    wire _3416;
    wire _4045;
    wire _4046;
    wire _4047;
    wire _4048;
    wire _4049;
    wire _4492;
    wire _3417;
    wire _4050;
    wire _4051;
    wire _4052;
    wire _4053;
    wire _4054;
    wire _4491;
    wire _3418;
    wire _4055;
    wire _4056;
    wire _4057;
    wire _4058;
    wire _4059;
    wire _4490;
    wire _3419;
    wire _4060;
    wire _4061;
    wire _4062;
    wire _4063;
    wire _4064;
    wire _4489;
    wire _3420;
    wire _4065;
    wire _4066;
    wire _4067;
    wire _4068;
    wire _4069;
    wire _4488;
    wire _3421;
    wire _4070;
    wire _4071;
    wire _4072;
    wire _4073;
    wire _4074;
    wire _4487;
    wire _3422;
    wire _4075;
    wire _4076;
    wire _4077;
    wire _4078;
    wire _4079;
    wire _4486;
    wire _3423;
    wire _4080;
    wire _4081;
    wire _4082;
    wire _4083;
    wire _4084;
    wire _4485;
    wire _3424;
    wire _4085;
    wire _4086;
    wire _4087;
    wire _4088;
    wire _4089;
    wire _4484;
    wire _3425;
    wire _4090;
    wire _4091;
    wire _4092;
    wire _4093;
    wire _4094;
    wire _4483;
    wire _3426;
    wire _4095;
    wire _4096;
    wire _4097;
    wire _4098;
    wire _4099;
    wire _4482;
    wire _3427;
    wire _4100;
    wire _4101;
    wire _4102;
    wire _4103;
    wire _4104;
    wire _4481;
    wire _3428;
    wire _4105;
    wire _4106;
    wire _4107;
    wire _4108;
    wire _4109;
    wire _4480;
    wire _3429;
    wire _4110;
    wire _4111;
    wire _4112;
    wire _4113;
    wire _4114;
    wire _4479;
    wire _3430;
    wire _4115;
    wire _4116;
    wire _4117;
    wire _4118;
    wire _4119;
    wire _4478;
    wire _3431;
    wire _4120;
    wire _4121;
    wire _4122;
    wire _4123;
    wire _4124;
    wire _4477;
    wire _3432;
    wire _4125;
    wire [31:0] _38 = 32'b11111111111111111111111111111111;
    wire _4126;
    wire _4127;
    wire _4128;
    wire _4129;
    wire _4476;
    wire _3433;
    wire [31:0] _3434;
    wire _4529;
    wire [31:0] _4530;
    wire [31:0] _3399;
    reg [31:0] _3401;
    wire _4910;
    wire _4911;
    wire _4912;
    wire _4913;
    wire _4914;
    wire _4915;
    wire _4916;
    wire _4917;
    wire _4918;
    wire _4919;
    wire _4920;
    wire _4921;
    wire _4922;
    wire _4923;
    wire _4924;
    wire _4925;
    wire _4926;
    wire _4927;
    wire _4928;
    wire _4929;
    wire _4930;
    wire _4931;
    wire _4932;
    wire _4933;
    wire _4934;
    wire _4935;
    wire _4936;
    wire _4937;
    wire _4938;
    wire _4939;
    wire _4940;
    wire _4941;
    wire _4942;
    wire _4943;
    wire _4944;
    wire _3946 = 1'b0;
    wire _4945;
    wire _4946;
    wire _3335;
    reg _3337;
    wire _3559;
    wire _3560;
    wire _3561;
    wire _4857;
    wire _4858;
    wire _3741 = 1'b1;
    wire _3744;
    wire _3745;
    wire _4859;
    wire _3749;
    wire _3750;
    wire _3751;
    wire _4860;
    wire _3753;
    wire _3754;
    wire _3755;
    wire _4861;
    wire _3759;
    wire _4862;
    wire _3775;
    wire _4863;
    wire _3790;
    wire _4864;
    wire _3809;
    wire _4865;
    wire _4866;
    wire _4867;
    wire _4868;
    wire _4869;
    wire _4870;
    wire _4871;
    wire _3347;
    reg _3349;
    wire [31:0] _4975;
    wire [31:0] _2673 = 32'b00000000000000000000000000000000;
    wire _4976;
    wire [31:0] _4977;
    wire [31:0] _2674;
    reg [31:0] _3070;
    reg [31:0] _3246;
    wire [31:0] _3686 = 32'b00000000000000000000000000000000;
    wire [5:0] _3687 = 6'b000000;
    wire _3688;
    wire _3689;
    wire [31:0] _3690;
    wire [4:0] _3806;
    wire [4:0] _3839 = 5'b00100;
    wire [4:0] _3840;
    wire [4:0] _3815 = 5'b00001;
    wire [4:0] _3816;
    wire [4:0] _3866 = 5'b00100;
    wire _3867;
    wire _3868;
    wire [4:0] _4561;
    wire [4:0] _4562;
    wire [4:0] _4131 = 5'b00000;
    wire _4563;
    wire [4:0] _4564;
    wire _4565;
    wire [4:0] _4566;
    wire _4567;
    wire [4:0] _4568;
    wire [4:0] _3387;
    reg [4:0] _3389;
    wire _3870;
    wire [31:0] _5003;
    wire [31:0] _3877;
    wire _2647 = 1'b0;
    wire _2645 = 1'b0;
    wire _3939 = 1'b1;
    wire _3942 = 1'b0;
    wire _5139;
    wire _3876 = 1'b1;
    wire _4152;
    wire _4153;
    wire _4154;
    wire _4155;
    wire _3532;
    wire _5140;
    wire _2646;
    reg _2648;
    wire _3888;
    wire [31:0] _5004;
    wire _3889;
    wire _3890;
    wire [31:0] _5005;
    wire [31:0] _3917;
    wire _2643 = 1'b0;
    wire _2641 = 1'b0;
    wire _3940 = 1'b1;
    wire _3943 = 1'b0;
    wire _5141;
    wire _3916 = 1'b1;
    wire _4148;
    wire _4149;
    wire _4150;
    wire _4151;
    wire _3533;
    wire _5142;
    wire _2642;
    reg _2644;
    wire _3935;
    wire [31:0] _5006;
    wire [31:0] _5007;
    wire _5008;
    wire [31:0] _5009;
    wire _5010;
    wire [31:0] _5011;
    wire _5012;
    wire [31:0] _5013;
    wire _5014;
    wire [31:0] _5015;
    wire [31:0] _2662;
    reg [31:0] _2664;
    wire _3248;
    wire _3259;
    wire _3279;
    wire _3262;
    wire _3273;
    wire _3282;
    wire _3276;
    wire _3278;
    wire _3284;
    wire _3286;
    wire _3287;
    wire _4144;
    wire _3813;
    wire _4145;
    wire gnd = 1'b0;
    wire _4146;
    wire _4147;
    wire _3534;
    wire _5138;
    wire _2650;
    reg _2652;
    wire _3948;
    wire _5176;
    wire _5177;
    wire _5178;
    wire _5179;
    wire _5180;
    wire _5181;
    wire _2626;
    reg _2628;
    wire _3651;
    wire _3652;
    wire _3653;
    wire vdd = 1'b1;
    wire _3654;
    wire _5156;
    wire _5157;
    wire _5158;
    wire _5159;
    wire _2634;
    reg _2636;
    wire _3936;
    wire _3937;
    wire [2:0] _5240;
    wire [2:0] _2598 = 3'b111;
    wire _5241;
    wire [2:0] _5242;
    wire [2:0] _2599 = 3'b110;
    wire _5243;
    wire [2:0] _5244;
    wire [2:0] _2600 = 3'b101;
    wire _5245;
    wire [2:0] _5246;
    wire [2:0] _2601 = 3'b100;
    wire _5247;
    wire [2:0] _5248;
    wire [2:0] _2602 = 3'b011;
    wire _5249;
    wire [2:0] _5250;
    wire [2:0] _2603 = 3'b010;
    wire _5251;
    wire [2:0] _5252;
    wire [2:0] _2605 = 3'b000;
    wire _5253;
    wire [2:0] _5254;
    wire [2:0] _2606;
    reg [2:0] _2608;
    wire _4848;
    wire _4849;
    wire _3355;
    reg _3357;
    wire _5255;
    wire [31:0] _5256;

    /* logic */
    assign _5296 = _2598 == _2608;
    assign _5444 = _5296 ? _5295 : _5275;
    assign _5317 = _2599 == _2608;
    assign _5445 = _5317 ? _5316 : _5444;
    assign _5338 = _2600 == _2608;
    assign _5446 = _5338 ? _5337 : _5445;
    assign _5359 = _2601 == _2608;
    assign _5447 = _5359 ? _5358 : _5446;
    assign _5380 = _2602 == _2608;
    assign _5448 = _5380 ? _5379 : _5447;
    assign _5401 = _2603 == _2608;
    assign _5449 = _5401 ? _5400 : _5448;
    assign _5422 = _2605 == _2608;
    assign _5450 = _5422 ? _5421 : _5449;
    assign _5443 = _2604 == _2608;
    assign ascii_state_0 = _5443 ? _5442 : _5450;
    assign _3664 = ~ _3531;
    assign _3665 = _3401 & _3664;
    assign _5190 = _3667 ? _3665 : _2616;
    assign _5191 = _3671 ? _2616 : _5190;
    assign _5192 = _3357 ? _2616 : _5191;
    assign _5193 = _3349 ? _2616 : _5192;
    assign _5194 = _3745 ? _3743 : _2616;
    assign _5195 = _3751 ? _2616 : _5194;
    assign _5196 = _3755 ? _2616 : _5195;
    assign _5197 = _3759 ? _2616 : _5196;
    assign _5198 = _3775 ? _2616 : _5197;
    assign _5199 = _3790 ? _2616 : _5198;
    assign _5200 = _2608 == _2603;
    assign _5201 = _5200 ? _5199 : _2616;
    assign _5202 = _2608 == _2605;
    assign _5203 = _5202 ? _5193 : _5201;
    assign _2614 = _5203;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2616 <= _2613;
        else
            _2616 <= _2614;
    end
    assign _5182 = _3875 ? _3872 : _3947;
    assign _5183 = _3890 ? _5182 : _3947;
    assign _5184 = _3915 ? _3891 : _3947;
    assign _5185 = _3937 ? _5184 : _3947;
    assign _5186 = _2608 == _2598;
    assign _5187 = _5186 ? _5185 : _3947;
    assign _5188 = _2608 == _2599;
    assign _5189 = _5188 ? _5183 : _5187;
    assign _2618 = _5189;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2620 <= _2617;
        else
            _2620 <= _2618;
    end
    assign _2622 = _2628;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2624 <= _2621;
        else
            _2624 <= _2622;
    end
    assign _3884 = _3883 ? _3882 : _3880;
    assign _3881 = instr[16:16];
    assign _3883 = instr[15:15];
    assign _3885 = _3883 | _3881;
    assign _3886 = _3885 ? _3884 : _3878;
    assign _5143 = _3888 ? _3886 : _2640;
    assign _5144 = _3890 ? _5143 : _2640;
    assign _3931 = _3930 ? _3927 : _3923;
    assign _3924 = instr[14:14];
    assign _3925 = instr[11:11];
    assign _3926 = _3925 | _3924;
    assign _3928 = instr[13:13];
    assign _3929 = instr[10:10];
    assign _3930 = _3929 | _3928;
    assign _3932 = _3930 | _3926;
    assign _3933 = _3932 ? _3931 : _3921;
    assign _5145 = _3935 ? _3933 : _2640;
    assign _5146 = _3937 ? _5145 : _2640;
    assign _5147 = _2608 == _2598;
    assign _5148 = _5147 ? _5146 : _2640;
    assign _5149 = _2608 == _2599;
    assign _5150 = _5149 ? _5144 : _5148;
    assign _5151 = _2608 == _2605;
    assign _5152 = _5151 ? _3677 : _5150;
    assign _2638 = _5152;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2640 <= _2637;
        else
            _2640 <= _2638;
    end
    assign _5034 = _2608 == _2604;
    assign _5035 = _5034 ? vdd : _4132;
    assign _2654 = _5035;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2656 <= _2653;
        else
            _2656 <= _2654;
    end
    assign _4758 = _3401[0:0];
    assign _4759 = _3401[1:1];
    assign _4760 = _3401[2:2];
    assign _4761 = _3401[3:3];
    assign _4762 = _3401[4:4];
    assign _4763 = _3401[5:5];
    assign _4764 = _3401[6:6];
    assign _4765 = _3401[7:7];
    assign _4766 = _3401[8:8];
    assign _4767 = _3401[9:9];
    assign _4768 = _3401[10:10];
    assign _4769 = _3401[11:11];
    assign _4770 = _3401[12:12];
    assign _4771 = _3401[13:13];
    assign _4772 = _3401[14:14];
    assign _4773 = _3401[15:15];
    assign _4774 = _3401[16:16];
    assign _4775 = _3401[17:17];
    assign _4776 = _3401[18:18];
    assign _4777 = _3401[19:19];
    assign _4778 = _3401[20:20];
    assign _4779 = _3401[21:21];
    assign _4780 = _3401[22:22];
    assign _4781 = _3401[23:23];
    assign _4782 = _3401[24:24];
    assign _4783 = _3401[25:25];
    assign _4784 = _3401[26:26];
    assign _4785 = _3401[27:27];
    assign _4786 = _3401[28:28];
    assign _4787 = _3401[29:29];
    assign _4788 = _3401[30:30];
    assign _4789 = _3401[31:31];
    assign _4790 = _4789 | _4788;
    assign _4791 = _4790 | _4787;
    assign _4792 = _4791 | _4786;
    assign _4793 = _4792 | _4785;
    assign _4794 = _4793 | _4784;
    assign _4795 = _4794 | _4783;
    assign _4796 = _4795 | _4782;
    assign _4797 = _4796 | _4781;
    assign _4798 = _4797 | _4780;
    assign _4799 = _4798 | _4779;
    assign _4800 = _4799 | _4778;
    assign _4801 = _4800 | _4777;
    assign _4802 = _4801 | _4776;
    assign _4803 = _4802 | _4775;
    assign _4804 = _4803 | _4774;
    assign _4805 = _4804 | _4773;
    assign _4806 = _4805 | _4772;
    assign _4807 = _4806 | _4771;
    assign _4808 = _4807 | _4770;
    assign _4809 = _4808 | _4769;
    assign _4810 = _4809 | _4768;
    assign _4811 = _4810 | _4767;
    assign _4812 = _4811 | _4766;
    assign _4813 = _4812 | _4765;
    assign _4814 = _4813 | _4764;
    assign _4815 = _4814 | _4763;
    assign _4816 = _4815 | _4762;
    assign _4817 = _4816 | _4761;
    assign _4818 = _4817 | _4760;
    assign _4819 = _4818 | _4759;
    assign _4820 = _4819 | _4758;
    assign _4821 = _4820 ? _3557 : _3660;
    assign _4822 = _3561 ? _4821 : _3660;
    assign _4823 = _3654 ? _3660 : _4822;
    assign _4824 = pcpi_int_ready ? pcpi_int_wr : _3357;
    assign _4825 = vdd ? _4824 : _3357;
    assign _4826 = vdd ? _4825 : _3357;
    assign _4827 = _3703 ? _3700 : _3357;
    assign _4828 = _3739 ? _3737 : _4827;
    assign _4829 = _3745 ? _3740 : _4828;
    assign _4830 = _3751 ? _3746 : _4829;
    assign _4831 = _3755 ? _3752 : _4830;
    assign _4832 = _3759 ? _3357 : _4831;
    assign _4833 = _3775 ? _3760 : _4832;
    assign _4834 = _3790 ? _4826 : _4833;
    assign _4835 = pcpi_int_ready ? pcpi_int_wr : _3357;
    assign _4836 = _3805 ? _4835 : _3357;
    assign _4837 = _3813 ? _3287 : _3808;
    assign _4838 = _2608 == _2598;
    assign _4839 = _4838 ? _3938 : _3357;
    assign _4840 = _2608 == _2600;
    assign _4841 = _4840 ? _3871 : _4839;
    assign _4842 = _2608 == _2601;
    assign _4843 = _4842 ? _4837 : _4841;
    assign _4844 = _2608 == _2602;
    assign _4845 = _4844 ? _4836 : _4843;
    assign _4846 = _2608 == _2603;
    assign _4847 = _4846 ? _4834 : _4845;
    assign _5204 = _3548 ? _2608 : _2603;
    assign _5205 = _2628 ? _5204 : _2608;
    assign _5206 = _3561 ? _2608 : _5205;
    assign _5207 = _3654 ? _2608 : _5206;
    assign _5208 = _3785 ? _2605 : _2604;
    assign _5209 = _3329 ? _5208 : _2608;
    assign _5210 = pcpi_int_ready ? _2605 : _5209;
    assign _5211 = vdd ? _5210 : _2602;
    assign _5212 = _3780 ? _2605 : _2604;
    assign _5213 = vdd ? _5211 : _5212;
    assign _5214 = _3691 ? _2600 : _2601;
    assign _5215 = _3693 ? _2599 : _5214;
    assign _5216 = vdd ? _5215 : _2602;
    assign _5217 = _3695 ? _2601 : _5216;
    assign _5218 = _3697 ? _2600 : _5217;
    assign _5219 = _3699 ? _2598 : _5218;
    assign _5220 = _3703 ? _2605 : _5219;
    assign _5221 = _3739 ? _2605 : _5220;
    assign _5222 = _3745 ? _2605 : _5221;
    assign _5223 = _3751 ? _2605 : _5222;
    assign _5224 = _3755 ? _2605 : _5223;
    assign _5225 = _3759 ? _2601 : _5224;
    assign _5226 = _3775 ? _2605 : _5225;
    assign _5227 = _3790 ? _5213 : _5226;
    assign _5228 = _3800 ? _2605 : _2604;
    assign _5229 = _3329 ? _5228 : _2608;
    assign _5230 = pcpi_int_ready ? _2605 : _5229;
    assign _5231 = _3793 ? _2600 : _2601;
    assign _5232 = _3795 ? _2599 : _5231;
    assign _5233 = _3805 ? _5230 : _5232;
    assign _5234 = mem_done ? _2605 : _2608;
    assign _5235 = _3813 ? _5234 : _2605;
    assign _5236 = _3870 ? _2605 : _2608;
    assign _5237 = _3875 ? _2605 : _2608;
    assign _5238 = _3890 ? _5237 : _2608;
    assign _5239 = _3915 ? _2605 : _2608;
    assign _3539 = instr[43:43];
    assign _3540 = ~ _3539;
    assign _3541 = instr[3:3];
    assign _3542 = ~ _3541;
    assign _3543 = _3542 & _3540;
    assign _5153 = _3548 ? _2636 : _3543;
    assign _5154 = _2628 ? _5153 : _2636;
    assign _5155 = _3561 ? _2636 : _5154;
    assign _3582 = _3393[0:0];
    assign _3583 = _3393[1:1];
    assign _3584 = _3583 | _3582;
    assign _3587 = _3586[0:0];
    assign _3588 = _3586[1:1];
    assign _3589 = _3586[2:2];
    assign _3590 = _3586[3:3];
    assign _3591 = _3586[4:4];
    assign _3592 = _3586[5:5];
    assign _3593 = _3586[6:6];
    assign _3594 = _3586[7:7];
    assign _3595 = _3586[8:8];
    assign _3596 = _3586[9:9];
    assign _3597 = _3586[10:10];
    assign _3598 = _3586[11:11];
    assign _3599 = _3586[12:12];
    assign _3600 = _3586[13:13];
    assign _3601 = _3586[14:14];
    assign _3602 = _3586[15:15];
    assign _3603 = _3586[16:16];
    assign _3604 = _3586[17:17];
    assign _3605 = _3586[18:18];
    assign _3606 = _3586[19:19];
    assign _3607 = _3586[20:20];
    assign _3608 = _3586[21:21];
    assign _3609 = _3586[22:22];
    assign _3610 = _3586[23:23];
    assign _3611 = _3586[24:24];
    assign _3612 = _3586[25:25];
    assign _3613 = _3586[26:26];
    assign _3614 = _3586[27:27];
    assign _3615 = _3586[28:28];
    assign _3616 = _3586[29:29];
    assign _3617 = _3586[30:30];
    assign _3585 = ~ _3531;
    assign _3586 = _3401 & _3585;
    assign _3618 = _3586[31:31];
    assign _3619 = _3618 | _3617;
    assign _3620 = _3619 | _3616;
    assign _3621 = _3620 | _3615;
    assign _3622 = _3621 | _3614;
    assign _3623 = _3622 | _3613;
    assign _3624 = _3623 | _3612;
    assign _3625 = _3624 | _3611;
    assign _3626 = _3625 | _3610;
    assign _3627 = _3626 | _3609;
    assign _3628 = _3627 | _3608;
    assign _3629 = _3628 | _3607;
    assign _3630 = _3629 | _3606;
    assign _3631 = _3630 | _3605;
    assign _3632 = _3631 | _3604;
    assign _3633 = _3632 | _3603;
    assign _3634 = _3633 | _3602;
    assign _3635 = _3634 | _3601;
    assign _3636 = _3635 | _3600;
    assign _3637 = _3636 | _3599;
    assign _3638 = _3637 | _3598;
    assign _3639 = _3638 | _3597;
    assign _3640 = _3639 | _3596;
    assign _3641 = _3640 | _3595;
    assign _3642 = _3641 | _3594;
    assign _3643 = _3642 | _3593;
    assign _3644 = _3643 | _3592;
    assign _3645 = _3644 | _3591;
    assign _3646 = _3645 | _3590;
    assign _3647 = _3646 | _3589;
    assign _3648 = _3647 | _3588;
    assign _3649 = _3648 | _3587;
    assign _3650 = ~ _3397;
    assign _5170 = _3287 ? _3811 : _3948;
    assign _5171 = _3813 ? _5170 : _3948;
    assign _3874 = ~ _2636;
    assign _3875 = _3874 & mem_done;
    assign _5172 = _3875 ? _3873 : _3948;
    assign _5173 = _3890 ? _5172 : _3948;
    assign _5174 = _3915 ? _3892 : _3948;
    assign _5175 = _3937 ? _5174 : _3948;
    assign _5039 = _3401[0:0];
    assign _5040 = _3401[1:1];
    assign _5041 = _3401[2:2];
    assign _5042 = _3401[3:3];
    assign _5043 = _3401[4:4];
    assign _5044 = _3401[5:5];
    assign _5045 = _3401[6:6];
    assign _5046 = _3401[7:7];
    assign _5047 = _3401[8:8];
    assign _5048 = _3401[9:9];
    assign _5049 = _3401[10:10];
    assign _5050 = _3401[11:11];
    assign _5051 = _3401[12:12];
    assign _5052 = _3401[13:13];
    assign _5053 = _3401[14:14];
    assign _5054 = _3401[15:15];
    assign _5055 = _3401[16:16];
    assign _5056 = _3401[17:17];
    assign _5057 = _3401[18:18];
    assign _5058 = _3401[19:19];
    assign _5059 = _3401[20:20];
    assign _5060 = _3401[21:21];
    assign _5061 = _3401[22:22];
    assign _5062 = _3401[23:23];
    assign _5063 = _3401[24:24];
    assign _5064 = _3401[25:25];
    assign _5065 = _3401[26:26];
    assign _5066 = _3401[27:27];
    assign _5067 = _3401[28:28];
    assign _5068 = _3401[29:29];
    assign _5069 = _3401[30:30];
    assign _5070 = _3401[31:31];
    assign _5071 = _5070 | _5069;
    assign _5072 = _5071 | _5068;
    assign _5073 = _5072 | _5067;
    assign _5074 = _5073 | _5066;
    assign _5075 = _5074 | _5065;
    assign _5076 = _5075 | _5064;
    assign _5077 = _5076 | _5063;
    assign _5078 = _5077 | _5062;
    assign _5079 = _5078 | _5061;
    assign _5080 = _5079 | _5060;
    assign _5081 = _5080 | _5059;
    assign _5082 = _5081 | _5058;
    assign _5083 = _5082 | _5057;
    assign _5084 = _5083 | _5056;
    assign _5085 = _5084 | _5055;
    assign _5086 = _5085 | _5054;
    assign _5087 = _5086 | _5053;
    assign _5088 = _5087 | _5052;
    assign _5089 = _5088 | _5051;
    assign _5090 = _5089 | _5050;
    assign _5091 = _5090 | _5049;
    assign _5092 = _5091 | _5048;
    assign _5093 = _5092 | _5047;
    assign _5094 = _5093 | _5046;
    assign _5095 = _5094 | _5045;
    assign _5096 = _5095 | _5044;
    assign _5097 = _5096 | _5043;
    assign _5098 = _5097 | _5042;
    assign _5099 = _5098 | _5041;
    assign _5100 = _5099 | _5040;
    assign _5101 = _5100 | _5039;
    assign _5102 = _5101 ? _3554 : _5038;
    assign _5103 = _3548 ? _3547 : _3544;
    assign _3678 = ~ _3337;
    assign _3679 = ~ _2628;
    assign _3680 = _3679 & _3678;
    assign _5036 = _3671 ? _3668 : _3680;
    assign _5037 = _3357 ? _3680 : _5036;
    assign _5038 = _3349 ? _3680 : _5037;
    assign _5104 = _2628 ? _5103 : _5038;
    assign _5105 = _3561 ? _5102 : _5104;
    assign _5106 = _3654 ? _5038 : _5105;
    assign _5107 = pcpi_int_ready ? _3787 : _2652;
    assign _5108 = vdd ? _5107 : _2652;
    assign _5109 = vdd ? _5108 : _2652;
    assign _3691 = is[5:5];
    assign _5110 = _3691 ? _2652 : _2636;
    assign _3693 = is[4:4];
    assign _5111 = _3693 ? _3692 : _5110;
    assign _5112 = vdd ? _5111 : _2652;
    assign _5113 = _3695 ? _2636 : _5112;
    assign _5114 = _3697 ? _2652 : _5113;
    assign _5115 = _3699 ? _3698 : _5114;
    assign _5116 = _3703 ? _2652 : _5115;
    assign _5117 = _3739 ? _2652 : _5116;
    assign _5118 = _3745 ? _2652 : _5117;
    assign _5119 = _3751 ? _2652 : _5118;
    assign _5120 = _3755 ? _2652 : _5119;
    assign _5121 = _3759 ? _2636 : _5120;
    assign _5122 = _3775 ? _2652 : _5121;
    assign _5123 = _3790 ? _5109 : _5122;
    assign _5124 = pcpi_int_ready ? _3802 : _2652;
    assign _3793 = is[5:5];
    assign _5125 = _3793 ? _2652 : _2636;
    assign _3795 = is[4:4];
    assign _5126 = _3795 ? _3794 : _5125;
    assign _5127 = _3805 ? _5124 : _5126;
    assign _5128 = _3870 ? _2636 : _2652;
    assign _5129 = _2608 == _2600;
    assign _5130 = _5129 ? _5128 : _2652;
    assign _5131 = _2608 == _2602;
    assign _5132 = _5131 ? _5127 : _5130;
    assign _5133 = _2608 == _2603;
    assign _5134 = _5133 ? _5123 : _5132;
    assign _5135 = _2608 == _2605;
    assign _5136 = _5135 ? _5106 : _5134;
    assign _5137 = mem_done ? _3944 : _5136;
    assign _3277 = _2664 == _2660;
    assign _3274 = _2664 == _2660;
    assign _3275 = ~ _3274;
    assign _3283 = _3278 ? _3277 : _3275;
    assign _3263 = _2660[30:0];
    assign _3264 = _2660[31:31];
    assign _3265 = ~ _3264;
    assign _3266 = { _3265, _3263 };
    assign _3267 = _2664[30:0];
    assign _3268 = _2664[31:31];
    assign _3269 = ~ _3268;
    assign _3270 = { _3269, _3267 };
    assign _3271 = _3270 < _3266;
    assign _3272 = ~ _3271;
    assign _3260 = _2664 < _2660;
    assign _3261 = ~ _3260;
    assign _3281 = _3273 ? _3272 : _3261;
    assign _3285 = _3284 ? _3283 : _3281;
    assign _3250 = _2660[30:0];
    assign _3251 = _2660[31:31];
    assign _3252 = ~ _3251;
    assign _3253 = { _3252, _3250 };
    assign _3254 = _2664[30:0];
    assign _3255 = _2664[31:31];
    assign _3256 = ~ _3255;
    assign _3257 = { _3256, _3254 };
    assign _3258 = _3257 < _3253;
    assign _4993 = vdd ? _3685 : _3792;
    assign _3757 = instr[0:0];
    assign _3758 = _3757 ? _3756 : _3375;
    assign _4994 = _3703 ? _3792 : _3685;
    assign _4995 = _3739 ? _3792 : _4994;
    assign _4996 = _3745 ? _3792 : _4995;
    assign _4997 = _3751 ? _3792 : _4996;
    assign _4998 = _3755 ? _3792 : _4997;
    assign _4999 = _3759 ? _3758 : _4998;
    assign _5000 = _3775 ? _3792 : _4999;
    assign _5001 = _3790 ? _4993 : _5000;
    assign _3857 = _2664[27:0];
    assign _3858 = { _3857, _3856 };
    assign _3850 = _2664[31:4];
    assign _3852 = { _3851, _3850 };
    assign _3862 = _3861 ? _3858 : _3852;
    assign _3841 = _2664[31:4];
    assign _3842 = _2664[31:31];
    assign _3843 = { _3842, _3842 };
    assign _3844 = { _3843, _3843 };
    assign _3846 = { _3844, _3841 };
    assign _3853 = instr[33:33];
    assign _3854 = instr[25:25];
    assign _3855 = _3854 | _3853;
    assign _3859 = instr[29:29];
    assign _3860 = instr[24:24];
    assign _3861 = _3860 | _3859;
    assign _3863 = _3861 | _3855;
    assign _3864 = _3863 ? _3862 : _3846;
    assign _3830 = _2664[30:0];
    assign _3831 = { _3830, _3829 };
    assign _3823 = _2664[31:1];
    assign _3825 = { _3824, _3823 };
    assign _3835 = _3834 ? _3831 : _3825;
    assign _3817 = _2664[31:1];
    assign _3818 = _2664[31:31];
    assign _3819 = { _3818, _3817 };
    assign _3826 = instr[33:33];
    assign _3827 = instr[25:25];
    assign _3828 = _3827 | _3826;
    assign _3832 = instr[29:29];
    assign _3833 = instr[24:24];
    assign _3834 = _3833 | _3832;
    assign _3836 = _3834 | _3828;
    assign _3837 = _3836 ? _3835 : _3819;
    assign _5002 = _3868 ? _3864 : _3837;
    assign _3788 = _3690[4:0];
    assign _4547 = vdd ? _3788 : _4131;
    assign _4548 = vdd ? _4547 : _4131;
    assign _3696 = decoded_rs2[4:0];
    assign _3694 = _3690[4:0];
    assign _4549 = vdd ? _3694 : _4131;
    assign _4550 = _3695 ? _4131 : _4549;
    assign _4551 = _3697 ? _3696 : _4550;
    assign _4552 = _3699 ? _4131 : _4551;
    assign _4553 = _3703 ? _4131 : _4552;
    assign _4554 = _3739 ? _4131 : _4553;
    assign _4555 = _3745 ? _4131 : _4554;
    assign _4556 = _3751 ? _4131 : _4555;
    assign _4557 = _3755 ? _4131 : _4556;
    assign _4558 = _3759 ? _4131 : _4557;
    assign _4559 = _3775 ? _4131 : _4558;
    assign _4560 = _3790 ? _4548 : _4559;
    assign _3066 = _3065[0:0];
    assign _3067 = _2675 & _3066;
    assign _3674 = _3375 + _3673;
    assign _4968 = vdd ? _3674 : _2673;
    assign _3672 = _3353 ? _3381 : _3385;
    assign _4969 = vdd ? _3672 : _2673;
    assign _3556 = _3377 + _3555;
    assign _4670 = _3401[0:0];
    assign _4671 = _3401[1:1];
    assign _4672 = _3401[2:2];
    assign _4673 = _3401[3:3];
    assign _4674 = _3401[4:4];
    assign _4675 = _3401[5:5];
    assign _4676 = _3401[6:6];
    assign _4677 = _3401[7:7];
    assign _4678 = _3401[8:8];
    assign _4679 = _3401[9:9];
    assign _4680 = _3401[10:10];
    assign _4681 = _3401[11:11];
    assign _4682 = _3401[12:12];
    assign _4683 = _3401[13:13];
    assign _4684 = _3401[14:14];
    assign _4685 = _3401[15:15];
    assign _4686 = _3401[16:16];
    assign _4687 = _3401[17:17];
    assign _4688 = _3401[18:18];
    assign _4689 = _3401[19:19];
    assign _4690 = _3401[20:20];
    assign _4691 = _3401[21:21];
    assign _4692 = _3401[22:22];
    assign _4693 = _3401[23:23];
    assign _4694 = _3401[24:24];
    assign _4695 = _3401[25:25];
    assign _4696 = _3401[26:26];
    assign _4697 = _3401[27:27];
    assign _4698 = _3401[28:28];
    assign _4699 = _3401[29:29];
    assign _4700 = _3401[30:30];
    assign _4701 = _3401[31:31];
    assign _4702 = _4701 | _4700;
    assign _4703 = _4702 | _4699;
    assign _4704 = _4703 | _4698;
    assign _4705 = _4704 | _4697;
    assign _4706 = _4705 | _4696;
    assign _4707 = _4706 | _4695;
    assign _4708 = _4707 | _4694;
    assign _4709 = _4708 | _4693;
    assign _4710 = _4709 | _4692;
    assign _4711 = _4710 | _4691;
    assign _4712 = _4711 | _4690;
    assign _4713 = _4712 | _4689;
    assign _4714 = _4713 | _4688;
    assign _4715 = _4714 | _4687;
    assign _4716 = _4715 | _4686;
    assign _4717 = _4716 | _4685;
    assign _4718 = _4717 | _4684;
    assign _4719 = _4718 | _4683;
    assign _4720 = _4719 | _4682;
    assign _4721 = _4720 | _4681;
    assign _4722 = _4721 | _4680;
    assign _4723 = _4722 | _4679;
    assign _4724 = _4723 | _4678;
    assign _4725 = _4724 | _4677;
    assign _4726 = _4725 | _4676;
    assign _4727 = _4726 | _4675;
    assign _4728 = _4727 | _4674;
    assign _4729 = _4728 | _4673;
    assign _4730 = _4729 | _4672;
    assign _4731 = _4730 | _4671;
    assign _4732 = _4731 | _4670;
    assign _4733 = _4732 ? _3556 : _3377;
    assign _3546 = _3377 + decoded_imm_uj;
    assign _3552 = _3377 + _3551;
    assign _4734 = _3548 ? _3546 : _3552;
    assign _3314 = _2664 + _2660;
    assign _3312 = _2664 - _2660;
    assign _3320 = _3315 ? _3314 : _3312;
    assign _3310 = { _3308, _3287 };
    assign _3297 = _2664 ^ _2660;
    assign _3318 = _3311 ? _3310 : _3297;
    assign _3322 = _3321 ? _3320 : _3318;
    assign _3293 = _2664 | _2660;
    assign _5016 = vdd ? _3690 : _3791;
    assign _5017 = vdd ? _5016 : _3791;
    assign _5018 = vdd ? _3690 : _3791;
    assign _3695 = is[3:3];
    assign _5019 = _3695 ? decoded_imm : _5018;
    assign _3697 = is[2:2];
    assign _5020 = _3697 ? _3791 : _5019;
    assign _3699 = is[1:1];
    assign _5021 = _3699 ? _3791 : _5020;
    assign _5022 = _3703 ? _3791 : _5021;
    assign _5023 = _3739 ? _3791 : _5022;
    assign _5024 = _3745 ? _3791 : _5023;
    assign _5025 = _3751 ? _3791 : _5024;
    assign _5026 = _3755 ? _3791 : _5025;
    assign _5027 = _3759 ? decoded_imm : _5026;
    assign _5028 = _3775 ? _3791 : _5027;
    assign _5029 = _3790 ? _5017 : _5028;
    assign _5030 = _2608 == _2602;
    assign _5031 = _5030 ? _3690 : _2660;
    assign _5032 = _2608 == _2603;
    assign _5033 = _5032 ? _5029 : _5031;
    assign _2658 = _5033;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2660 <= _2657;
        else
            _2660 <= _2658;
    end
    assign _3289 = _2664 & _2660;
    assign _3294 = instr[35:35];
    assign _3295 = instr[22:22];
    assign _3296 = _3295 | _3294;
    assign _3316 = _3296 ? _3293 : _3289;
    assign _3298 = instr[32:32];
    assign _3299 = instr[21:21];
    assign _3300 = _3299 | _3298;
    assign _3311 = is[13:13];
    assign _3319 = _3311 | _3300;
    assign _3313 = instr[28:28];
    assign _3315 = is[6:6];
    assign _3321 = _3315 | _3313;
    assign _3323 = _3321 | _3319;
    assign _3324 = _3323 ? _3322 : _3316;
    assign _3379 = _3324;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3381 <= _3378;
        else
            _3381 <= _3379;
    end
    assign _4569 = _3401[0:0];
    assign _4570 = _3401[1:1];
    assign _4571 = _3401[2:2];
    assign _4572 = _3401[3:3];
    assign _4573 = _3401[4:4];
    assign _4574 = _3401[5:5];
    assign _4575 = _3401[6:6];
    assign _4576 = _3401[7:7];
    assign _4577 = _3401[8:8];
    assign _4578 = _3401[9:9];
    assign _4579 = _3401[10:10];
    assign _4580 = _3401[11:11];
    assign _4581 = _3401[12:12];
    assign _4582 = _3401[13:13];
    assign _4583 = _3401[14:14];
    assign _4584 = _3401[15:15];
    assign _4585 = _3401[16:16];
    assign _4586 = _3401[17:17];
    assign _4587 = _3401[18:18];
    assign _4588 = _3401[19:19];
    assign _4589 = _3401[20:20];
    assign _4590 = _3401[21:21];
    assign _4591 = _3401[22:22];
    assign _4592 = _3401[23:23];
    assign _4593 = _3401[24:24];
    assign _4594 = _3401[25:25];
    assign _4595 = _3401[26:26];
    assign _4596 = _3401[27:27];
    assign _4597 = _3401[28:28];
    assign _4598 = _3401[29:29];
    assign _4599 = _3401[30:30];
    assign _4600 = _3401[31:31];
    assign _4601 = _4600 | _4599;
    assign _4602 = _4601 | _4598;
    assign _4603 = _4602 | _4597;
    assign _4604 = _4603 | _4596;
    assign _4605 = _4604 | _4595;
    assign _4606 = _4605 | _4594;
    assign _4607 = _4606 | _4593;
    assign _4608 = _4607 | _4592;
    assign _4609 = _4608 | _4591;
    assign _4610 = _4609 | _4590;
    assign _4611 = _4610 | _4589;
    assign _4612 = _4611 | _4588;
    assign _4613 = _4612 | _4587;
    assign _4614 = _4613 | _4586;
    assign _4615 = _4614 | _4585;
    assign _4616 = _4615 | _4584;
    assign _4617 = _4616 | _4583;
    assign _4618 = _4617 | _4582;
    assign _4619 = _4618 | _4581;
    assign _4620 = _4619 | _4580;
    assign _4621 = _4620 | _4579;
    assign _4622 = _4621 | _4578;
    assign _4623 = _4622 | _4577;
    assign _4624 = _4623 | _4576;
    assign _4625 = _4624 | _4575;
    assign _4626 = _4625 | _4574;
    assign _4627 = _4626 | _4573;
    assign _4628 = _4627 | _4572;
    assign _4629 = _4628 | _4571;
    assign _4630 = _4629 | _4570;
    assign _4631 = _4630 | _4569;
    assign _4632 = _4631 ? _3401 : _4130;
    assign _4633 = _3561 ? _4632 : _4130;
    assign _4634 = _3654 ? _4130 : _4633;
    assign _4635 = pcpi_int_ready ? pcpi_int_rd : _4130;
    assign _4636 = vdd ? _4635 : _4130;
    assign _4637 = vdd ? _4636 : _4130;
    assign _3767 = count_cycle[31:0];
    assign _3962 = count_cycle + _3961;
    assign _4872 = vdd ? _3962 : count_cycle;
    assign _3343 = _4872;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            count_cycle <= _3342;
        else
            count_cycle <= _3343;
    end
    assign _3765 = count_cycle[63:32];
    assign _3771 = _3768 ? _3767 : _3765;
    assign _3763 = _3341[31:0];
    assign _3550 = _3341 + _3549;
    assign _4873 = vdd ? _3550 : _3341;
    assign _4874 = _2628 ? _4873 : _3341;
    assign _4875 = _3561 ? _3341 : _4874;
    assign _4876 = _3654 ? _3341 : _4875;
    assign _4877 = _2608 == _2605;
    assign _4878 = _4877 ? _4876 : _3341;
    assign _3339 = _4878;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3341 <= _3338;
        else
            _3341 <= _3339;
    end
    assign _3761 = _3341[63:32];
    assign _3764 = instr[39:39];
    assign _3769 = _3764 ? _3763 : _3761;
    assign _3766 = instr[38:38];
    assign _3768 = instr[37:37];
    assign _3772 = _3768 | _3766;
    assign _3773 = _3772 ? _3771 : _3769;
    assign _4638 = _3703 ? _3538 : _4130;
    assign _4639 = _3739 ? _3531 : _4638;
    assign _4640 = _3745 ? _3247 : _4639;
    assign _4641 = _3751 ? _3247 : _4640;
    assign _4642 = _3755 ? _3247 : _4641;
    assign _4643 = _3759 ? _4130 : _4642;
    assign _4644 = _3775 ? _3773 : _4643;
    assign _4645 = _3790 ? _4637 : _4644;
    assign _4646 = pcpi_int_ready ? pcpi_int_rd : _4130;
    assign _4647 = _3805 ? _4646 : _4130;
    assign _4668 = _2608 == _2605;
    assign _4669 = _4668 ? _3377 : _3375;
    assign _3373 = _4669;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3375 <= _39;
        else
            _3375 <= _3373;
    end
    assign _3814 = _3375 + decoded_imm;
    assign _4648 = _3870 ? _2664 : _4130;
    assign _3902 = mem_rdata_word[15:0];
    assign _3903 = _3902[15:15];
    assign _3904 = { _3903, _3903 };
    assign _3905 = { _3904, _3904 };
    assign _3906 = { _3905, _3905 };
    assign _3907 = { _3906, _3906 };
    assign _3909 = { _3907, _3902 };
    assign _3910 = _3369 ? mem_rdata_word : _3909;
    assign _3893 = mem_rdata_word[7:0];
    assign _3894 = _3893[7:7];
    assign _3895 = { _3894, _3894 };
    assign _3896 = { _3895, _3895 };
    assign _3897 = { _3896, _3896 };
    assign _3898 = { _3897, _3897 };
    assign _3899 = { _3898, _3897 };
    assign _3901 = { _3899, _3893 };
    assign _3919 = instr[11:11];
    assign _4746 = _3935 ? _3919 : _3365;
    assign _4747 = _3937 ? _4746 : _3365;
    assign _4748 = _2608 == _2598;
    assign _4749 = _4748 ? _4747 : _3365;
    assign _4750 = _2608 == _2605;
    assign _4751 = _4750 ? _3656 : _4749;
    assign _3363 = _4751;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3365 <= _3362;
        else
            _3365 <= _3363;
    end
    assign _3920 = is[10:10];
    assign _4740 = _3935 ? _3920 : _3369;
    assign _4741 = _3937 ? _4740 : _3369;
    assign _4742 = _2608 == _2598;
    assign _4743 = _4742 ? _4741 : _3369;
    assign _4744 = _2608 == _2605;
    assign _4745 = _4744 ? _3657 : _4743;
    assign _3367 = _4745;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3369 <= _3366;
        else
            _3369 <= _3367;
    end
    assign _3911 = _3369 | _3365;
    assign _3912 = _3911 ? _3910 : _3901;
    assign _3914 = ~ _2636;
    assign _3915 = _3914 & mem_done;
    assign _4649 = _3915 ? _3912 : _4130;
    assign _4650 = _3937 ? _4649 : _4130;
    assign _4651 = _2608 == _2598;
    assign _4652 = _4651 ? _4650 : _4130;
    assign _4653 = _2608 == _2600;
    assign _4654 = _4653 ? _4648 : _4652;
    assign _4655 = _2608 == _2601;
    assign _4656 = _4655 ? _3814 : _4654;
    assign _4657 = _2608 == _2602;
    assign _4658 = _4657 ? _4647 : _4656;
    assign _4659 = _2608 == _2603;
    assign _4660 = _4659 ? _4645 : _4658;
    assign _4661 = _2608 == _2605;
    assign _4662 = _4661 ? _4634 : _4660;
    assign _3383 = _4662;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3385 <= _3382;
        else
            _3385 <= _3383;
    end
    assign _4850 = _3813 ? _3353 : _3807;
    assign _4851 = _2608 == _2601;
    assign _4852 = _4851 ? _4850 : _3353;
    assign _4853 = _2608 == _2605;
    assign _4854 = _4853 ? _3659 : _4852;
    assign _3351 = _4854;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3353 <= _3350;
        else
            _3353 <= _3351;
    end
    assign _3675 = _3353 ? _3381 : _3385;
    assign _3676 = _3357 ? _3675 : _3372;
    assign _4663 = _3671 ? _40 : _3372;
    assign _4664 = _3357 ? _3372 : _4663;
    assign _4665 = _3349 ? _3676 : _4664;
    assign _4666 = _2608 == _2605;
    assign _4667 = _4666 ? _4665 : _3376;
    assign _3377 = _4667;
    assign _4735 = _2628 ? _4734 : _3377;
    assign _4736 = _3561 ? _4733 : _4735;
    assign _4737 = _3654 ? _3377 : _4736;
    assign _4738 = _2608 == _2605;
    assign _4739 = _4738 ? _4737 : _3372;
    assign _3370 = _4739;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3372 <= _39;
        else
            _3372 <= _3370;
    end
    assign _4970 = vdd ? _3372 : _2673;
    assign _3662 = ~ _3531;
    assign _3663 = _3401 & _3662;
    assign _4971 = vdd ? _3663 : _2673;
    assign _4972 = _3667 ? _4971 : _2673;
    assign _4973 = _3671 ? _4970 : _4972;
    assign _4974 = _3357 ? _4969 : _4973;
    assign _3548 = instr[2:2];
    assign _4855 = _3548 ? _3545 : _3658;
    assign _4856 = _2628 ? _4855 : _3658;
    assign _3558 = instr[45:45];
    assign _4879 = _3401[0:0];
    assign _4880 = _3401[1:1];
    assign _4881 = _3401[2:2];
    assign _4882 = _3401[3:3];
    assign _4883 = _3401[4:4];
    assign _4884 = _3401[5:5];
    assign _4885 = _3401[6:6];
    assign _4886 = _3401[7:7];
    assign _4887 = _3401[8:8];
    assign _4888 = _3401[9:9];
    assign _4889 = _3401[10:10];
    assign _4890 = _3401[11:11];
    assign _4891 = _3401[12:12];
    assign _4892 = _3401[13:13];
    assign _4893 = _3401[14:14];
    assign _4894 = _3401[15:15];
    assign _4895 = _3401[16:16];
    assign _4896 = _3401[17:17];
    assign _4897 = _3401[18:18];
    assign _4898 = _3401[19:19];
    assign _4899 = _3401[20:20];
    assign _4900 = _3401[21:21];
    assign _4901 = _3401[22:22];
    assign _4902 = _3401[23:23];
    assign _4903 = _3401[24:24];
    assign _4904 = _3401[25:25];
    assign _4905 = _3401[26:26];
    assign _4906 = _3401[27:27];
    assign _4907 = _3401[28:28];
    assign _4908 = _3401[29:29];
    assign _4909 = _3401[30:30];
    assign _3705 = _3704[0:0];
    assign _4466 = vdd ? _3705 : _3437;
    assign _4467 = _3739 ? _4466 : _3437;
    assign _4468 = _3745 ? _3437 : _4467;
    assign _4469 = _3751 ? _3437 : _4468;
    assign _4470 = _3755 ? _3437 : _4469;
    assign _4471 = _3759 ? _3437 : _4470;
    assign _4472 = _3775 ? _3437 : _4471;
    assign _4473 = _3790 ? _3437 : _4472;
    assign _4474 = _2608 == _2603;
    assign _4475 = _4474 ? _4473 : _3437;
    assign _3435 = _4475;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3437 <= vdd;
        else
            _3437 <= _3435;
    end
    assign _3707 = _3704[2:2];
    assign _4446 = vdd ? _3707 : _3443;
    assign _4447 = _3739 ? _4446 : _3443;
    assign _4448 = _3745 ? _3443 : _4447;
    assign _4449 = _3751 ? _3443 : _4448;
    assign _4450 = _3755 ? _3443 : _4449;
    assign _4451 = _3759 ? _3443 : _4450;
    assign _4452 = _3775 ? _3443 : _4451;
    assign _4453 = _3790 ? _3443 : _4452;
    assign _4454 = _2608 == _2603;
    assign _4455 = _4454 ? _4453 : _3443;
    assign _3441 = _4455;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3443 <= vdd;
        else
            _3443 <= _3441;
    end
    assign _3708 = _3704[3:3];
    assign _4436 = vdd ? _3708 : _3446;
    assign _4437 = _3739 ? _4436 : _3446;
    assign _4438 = _3745 ? _3446 : _4437;
    assign _4439 = _3751 ? _3446 : _4438;
    assign _4440 = _3755 ? _3446 : _4439;
    assign _4441 = _3759 ? _3446 : _4440;
    assign _4442 = _3775 ? _3446 : _4441;
    assign _4443 = _3790 ? _3446 : _4442;
    assign _4444 = _2608 == _2603;
    assign _4445 = _4444 ? _4443 : _3446;
    assign _3444 = _4445;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3446 <= vdd;
        else
            _3446 <= _3444;
    end
    assign _3709 = _3704[4:4];
    assign _4426 = vdd ? _3709 : _3449;
    assign _4427 = _3739 ? _4426 : _3449;
    assign _4428 = _3745 ? _3449 : _4427;
    assign _4429 = _3751 ? _3449 : _4428;
    assign _4430 = _3755 ? _3449 : _4429;
    assign _4431 = _3759 ? _3449 : _4430;
    assign _4432 = _3775 ? _3449 : _4431;
    assign _4433 = _3790 ? _3449 : _4432;
    assign _4434 = _2608 == _2603;
    assign _4435 = _4434 ? _4433 : _3449;
    assign _3447 = _4435;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3449 <= vdd;
        else
            _3449 <= _3447;
    end
    assign _3710 = _3704[5:5];
    assign _4416 = vdd ? _3710 : _3452;
    assign _4417 = _3739 ? _4416 : _3452;
    assign _4418 = _3745 ? _3452 : _4417;
    assign _4419 = _3751 ? _3452 : _4418;
    assign _4420 = _3755 ? _3452 : _4419;
    assign _4421 = _3759 ? _3452 : _4420;
    assign _4422 = _3775 ? _3452 : _4421;
    assign _4423 = _3790 ? _3452 : _4422;
    assign _4424 = _2608 == _2603;
    assign _4425 = _4424 ? _4423 : _3452;
    assign _3450 = _4425;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3452 <= vdd;
        else
            _3452 <= _3450;
    end
    assign _3711 = _3704[6:6];
    assign _4406 = vdd ? _3711 : _3455;
    assign _4407 = _3739 ? _4406 : _3455;
    assign _4408 = _3745 ? _3455 : _4407;
    assign _4409 = _3751 ? _3455 : _4408;
    assign _4410 = _3755 ? _3455 : _4409;
    assign _4411 = _3759 ? _3455 : _4410;
    assign _4412 = _3775 ? _3455 : _4411;
    assign _4413 = _3790 ? _3455 : _4412;
    assign _4414 = _2608 == _2603;
    assign _4415 = _4414 ? _4413 : _3455;
    assign _3453 = _4415;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3455 <= vdd;
        else
            _3455 <= _3453;
    end
    assign _3712 = _3704[7:7];
    assign _4396 = vdd ? _3712 : _3458;
    assign _4397 = _3739 ? _4396 : _3458;
    assign _4398 = _3745 ? _3458 : _4397;
    assign _4399 = _3751 ? _3458 : _4398;
    assign _4400 = _3755 ? _3458 : _4399;
    assign _4401 = _3759 ? _3458 : _4400;
    assign _4402 = _3775 ? _3458 : _4401;
    assign _4403 = _3790 ? _3458 : _4402;
    assign _4404 = _2608 == _2603;
    assign _4405 = _4404 ? _4403 : _3458;
    assign _3456 = _4405;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3458 <= vdd;
        else
            _3458 <= _3456;
    end
    assign _3713 = _3704[8:8];
    assign _4386 = vdd ? _3713 : _3461;
    assign _4387 = _3739 ? _4386 : _3461;
    assign _4388 = _3745 ? _3461 : _4387;
    assign _4389 = _3751 ? _3461 : _4388;
    assign _4390 = _3755 ? _3461 : _4389;
    assign _4391 = _3759 ? _3461 : _4390;
    assign _4392 = _3775 ? _3461 : _4391;
    assign _4393 = _3790 ? _3461 : _4392;
    assign _4394 = _2608 == _2603;
    assign _4395 = _4394 ? _4393 : _3461;
    assign _3459 = _4395;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3461 <= vdd;
        else
            _3461 <= _3459;
    end
    assign _3714 = _3704[9:9];
    assign _4376 = vdd ? _3714 : _3464;
    assign _4377 = _3739 ? _4376 : _3464;
    assign _4378 = _3745 ? _3464 : _4377;
    assign _4379 = _3751 ? _3464 : _4378;
    assign _4380 = _3755 ? _3464 : _4379;
    assign _4381 = _3759 ? _3464 : _4380;
    assign _4382 = _3775 ? _3464 : _4381;
    assign _4383 = _3790 ? _3464 : _4382;
    assign _4384 = _2608 == _2603;
    assign _4385 = _4384 ? _4383 : _3464;
    assign _3462 = _4385;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3464 <= vdd;
        else
            _3464 <= _3462;
    end
    assign _3715 = _3704[10:10];
    assign _4366 = vdd ? _3715 : _3467;
    assign _4367 = _3739 ? _4366 : _3467;
    assign _4368 = _3745 ? _3467 : _4367;
    assign _4369 = _3751 ? _3467 : _4368;
    assign _4370 = _3755 ? _3467 : _4369;
    assign _4371 = _3759 ? _3467 : _4370;
    assign _4372 = _3775 ? _3467 : _4371;
    assign _4373 = _3790 ? _3467 : _4372;
    assign _4374 = _2608 == _2603;
    assign _4375 = _4374 ? _4373 : _3467;
    assign _3465 = _4375;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3467 <= vdd;
        else
            _3467 <= _3465;
    end
    assign _3716 = _3704[11:11];
    assign _4356 = vdd ? _3716 : _3470;
    assign _4357 = _3739 ? _4356 : _3470;
    assign _4358 = _3745 ? _3470 : _4357;
    assign _4359 = _3751 ? _3470 : _4358;
    assign _4360 = _3755 ? _3470 : _4359;
    assign _4361 = _3759 ? _3470 : _4360;
    assign _4362 = _3775 ? _3470 : _4361;
    assign _4363 = _3790 ? _3470 : _4362;
    assign _4364 = _2608 == _2603;
    assign _4365 = _4364 ? _4363 : _3470;
    assign _3468 = _4365;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3470 <= vdd;
        else
            _3470 <= _3468;
    end
    assign _3717 = _3704[12:12];
    assign _4346 = vdd ? _3717 : _3473;
    assign _4347 = _3739 ? _4346 : _3473;
    assign _4348 = _3745 ? _3473 : _4347;
    assign _4349 = _3751 ? _3473 : _4348;
    assign _4350 = _3755 ? _3473 : _4349;
    assign _4351 = _3759 ? _3473 : _4350;
    assign _4352 = _3775 ? _3473 : _4351;
    assign _4353 = _3790 ? _3473 : _4352;
    assign _4354 = _2608 == _2603;
    assign _4355 = _4354 ? _4353 : _3473;
    assign _3471 = _4355;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3473 <= vdd;
        else
            _3473 <= _3471;
    end
    assign _3718 = _3704[13:13];
    assign _4336 = vdd ? _3718 : _3476;
    assign _4337 = _3739 ? _4336 : _3476;
    assign _4338 = _3745 ? _3476 : _4337;
    assign _4339 = _3751 ? _3476 : _4338;
    assign _4340 = _3755 ? _3476 : _4339;
    assign _4341 = _3759 ? _3476 : _4340;
    assign _4342 = _3775 ? _3476 : _4341;
    assign _4343 = _3790 ? _3476 : _4342;
    assign _4344 = _2608 == _2603;
    assign _4345 = _4344 ? _4343 : _3476;
    assign _3474 = _4345;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3476 <= vdd;
        else
            _3476 <= _3474;
    end
    assign _3719 = _3704[14:14];
    assign _4326 = vdd ? _3719 : _3479;
    assign _4327 = _3739 ? _4326 : _3479;
    assign _4328 = _3745 ? _3479 : _4327;
    assign _4329 = _3751 ? _3479 : _4328;
    assign _4330 = _3755 ? _3479 : _4329;
    assign _4331 = _3759 ? _3479 : _4330;
    assign _4332 = _3775 ? _3479 : _4331;
    assign _4333 = _3790 ? _3479 : _4332;
    assign _4334 = _2608 == _2603;
    assign _4335 = _4334 ? _4333 : _3479;
    assign _3477 = _4335;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3479 <= vdd;
        else
            _3479 <= _3477;
    end
    assign _3720 = _3704[15:15];
    assign _4316 = vdd ? _3720 : _3482;
    assign _4317 = _3739 ? _4316 : _3482;
    assign _4318 = _3745 ? _3482 : _4317;
    assign _4319 = _3751 ? _3482 : _4318;
    assign _4320 = _3755 ? _3482 : _4319;
    assign _4321 = _3759 ? _3482 : _4320;
    assign _4322 = _3775 ? _3482 : _4321;
    assign _4323 = _3790 ? _3482 : _4322;
    assign _4324 = _2608 == _2603;
    assign _4325 = _4324 ? _4323 : _3482;
    assign _3480 = _4325;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3482 <= vdd;
        else
            _3482 <= _3480;
    end
    assign _3721 = _3704[16:16];
    assign _4306 = vdd ? _3721 : _3485;
    assign _4307 = _3739 ? _4306 : _3485;
    assign _4308 = _3745 ? _3485 : _4307;
    assign _4309 = _3751 ? _3485 : _4308;
    assign _4310 = _3755 ? _3485 : _4309;
    assign _4311 = _3759 ? _3485 : _4310;
    assign _4312 = _3775 ? _3485 : _4311;
    assign _4313 = _3790 ? _3485 : _4312;
    assign _4314 = _2608 == _2603;
    assign _4315 = _4314 ? _4313 : _3485;
    assign _3483 = _4315;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3485 <= vdd;
        else
            _3485 <= _3483;
    end
    assign _3722 = _3704[17:17];
    assign _4296 = vdd ? _3722 : _3488;
    assign _4297 = _3739 ? _4296 : _3488;
    assign _4298 = _3745 ? _3488 : _4297;
    assign _4299 = _3751 ? _3488 : _4298;
    assign _4300 = _3755 ? _3488 : _4299;
    assign _4301 = _3759 ? _3488 : _4300;
    assign _4302 = _3775 ? _3488 : _4301;
    assign _4303 = _3790 ? _3488 : _4302;
    assign _4304 = _2608 == _2603;
    assign _4305 = _4304 ? _4303 : _3488;
    assign _3486 = _4305;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3488 <= vdd;
        else
            _3488 <= _3486;
    end
    assign _3723 = _3704[18:18];
    assign _4286 = vdd ? _3723 : _3491;
    assign _4287 = _3739 ? _4286 : _3491;
    assign _4288 = _3745 ? _3491 : _4287;
    assign _4289 = _3751 ? _3491 : _4288;
    assign _4290 = _3755 ? _3491 : _4289;
    assign _4291 = _3759 ? _3491 : _4290;
    assign _4292 = _3775 ? _3491 : _4291;
    assign _4293 = _3790 ? _3491 : _4292;
    assign _4294 = _2608 == _2603;
    assign _4295 = _4294 ? _4293 : _3491;
    assign _3489 = _4295;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3491 <= vdd;
        else
            _3491 <= _3489;
    end
    assign _3724 = _3704[19:19];
    assign _4276 = vdd ? _3724 : _3494;
    assign _4277 = _3739 ? _4276 : _3494;
    assign _4278 = _3745 ? _3494 : _4277;
    assign _4279 = _3751 ? _3494 : _4278;
    assign _4280 = _3755 ? _3494 : _4279;
    assign _4281 = _3759 ? _3494 : _4280;
    assign _4282 = _3775 ? _3494 : _4281;
    assign _4283 = _3790 ? _3494 : _4282;
    assign _4284 = _2608 == _2603;
    assign _4285 = _4284 ? _4283 : _3494;
    assign _3492 = _4285;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3494 <= vdd;
        else
            _3494 <= _3492;
    end
    assign _3725 = _3704[20:20];
    assign _4266 = vdd ? _3725 : _3497;
    assign _4267 = _3739 ? _4266 : _3497;
    assign _4268 = _3745 ? _3497 : _4267;
    assign _4269 = _3751 ? _3497 : _4268;
    assign _4270 = _3755 ? _3497 : _4269;
    assign _4271 = _3759 ? _3497 : _4270;
    assign _4272 = _3775 ? _3497 : _4271;
    assign _4273 = _3790 ? _3497 : _4272;
    assign _4274 = _2608 == _2603;
    assign _4275 = _4274 ? _4273 : _3497;
    assign _3495 = _4275;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3497 <= vdd;
        else
            _3497 <= _3495;
    end
    assign _3726 = _3704[21:21];
    assign _4256 = vdd ? _3726 : _3500;
    assign _4257 = _3739 ? _4256 : _3500;
    assign _4258 = _3745 ? _3500 : _4257;
    assign _4259 = _3751 ? _3500 : _4258;
    assign _4260 = _3755 ? _3500 : _4259;
    assign _4261 = _3759 ? _3500 : _4260;
    assign _4262 = _3775 ? _3500 : _4261;
    assign _4263 = _3790 ? _3500 : _4262;
    assign _4264 = _2608 == _2603;
    assign _4265 = _4264 ? _4263 : _3500;
    assign _3498 = _4265;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3500 <= vdd;
        else
            _3500 <= _3498;
    end
    assign _3727 = _3704[22:22];
    assign _4246 = vdd ? _3727 : _3503;
    assign _4247 = _3739 ? _4246 : _3503;
    assign _4248 = _3745 ? _3503 : _4247;
    assign _4249 = _3751 ? _3503 : _4248;
    assign _4250 = _3755 ? _3503 : _4249;
    assign _4251 = _3759 ? _3503 : _4250;
    assign _4252 = _3775 ? _3503 : _4251;
    assign _4253 = _3790 ? _3503 : _4252;
    assign _4254 = _2608 == _2603;
    assign _4255 = _4254 ? _4253 : _3503;
    assign _3501 = _4255;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3503 <= vdd;
        else
            _3503 <= _3501;
    end
    assign _3728 = _3704[23:23];
    assign _4236 = vdd ? _3728 : _3506;
    assign _4237 = _3739 ? _4236 : _3506;
    assign _4238 = _3745 ? _3506 : _4237;
    assign _4239 = _3751 ? _3506 : _4238;
    assign _4240 = _3755 ? _3506 : _4239;
    assign _4241 = _3759 ? _3506 : _4240;
    assign _4242 = _3775 ? _3506 : _4241;
    assign _4243 = _3790 ? _3506 : _4242;
    assign _4244 = _2608 == _2603;
    assign _4245 = _4244 ? _4243 : _3506;
    assign _3504 = _4245;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3506 <= vdd;
        else
            _3506 <= _3504;
    end
    assign _3729 = _3704[24:24];
    assign _4226 = vdd ? _3729 : _3509;
    assign _4227 = _3739 ? _4226 : _3509;
    assign _4228 = _3745 ? _3509 : _4227;
    assign _4229 = _3751 ? _3509 : _4228;
    assign _4230 = _3755 ? _3509 : _4229;
    assign _4231 = _3759 ? _3509 : _4230;
    assign _4232 = _3775 ? _3509 : _4231;
    assign _4233 = _3790 ? _3509 : _4232;
    assign _4234 = _2608 == _2603;
    assign _4235 = _4234 ? _4233 : _3509;
    assign _3507 = _4235;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3509 <= vdd;
        else
            _3509 <= _3507;
    end
    assign _3730 = _3704[25:25];
    assign _4216 = vdd ? _3730 : _3512;
    assign _4217 = _3739 ? _4216 : _3512;
    assign _4218 = _3745 ? _3512 : _4217;
    assign _4219 = _3751 ? _3512 : _4218;
    assign _4220 = _3755 ? _3512 : _4219;
    assign _4221 = _3759 ? _3512 : _4220;
    assign _4222 = _3775 ? _3512 : _4221;
    assign _4223 = _3790 ? _3512 : _4222;
    assign _4224 = _2608 == _2603;
    assign _4225 = _4224 ? _4223 : _3512;
    assign _3510 = _4225;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3512 <= vdd;
        else
            _3512 <= _3510;
    end
    assign _3731 = _3704[26:26];
    assign _4206 = vdd ? _3731 : _3515;
    assign _4207 = _3739 ? _4206 : _3515;
    assign _4208 = _3745 ? _3515 : _4207;
    assign _4209 = _3751 ? _3515 : _4208;
    assign _4210 = _3755 ? _3515 : _4209;
    assign _4211 = _3759 ? _3515 : _4210;
    assign _4212 = _3775 ? _3515 : _4211;
    assign _4213 = _3790 ? _3515 : _4212;
    assign _4214 = _2608 == _2603;
    assign _4215 = _4214 ? _4213 : _3515;
    assign _3513 = _4215;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3515 <= vdd;
        else
            _3515 <= _3513;
    end
    assign _3732 = _3704[27:27];
    assign _4196 = vdd ? _3732 : _3518;
    assign _4197 = _3739 ? _4196 : _3518;
    assign _4198 = _3745 ? _3518 : _4197;
    assign _4199 = _3751 ? _3518 : _4198;
    assign _4200 = _3755 ? _3518 : _4199;
    assign _4201 = _3759 ? _3518 : _4200;
    assign _4202 = _3775 ? _3518 : _4201;
    assign _4203 = _3790 ? _3518 : _4202;
    assign _4204 = _2608 == _2603;
    assign _4205 = _4204 ? _4203 : _3518;
    assign _3516 = _4205;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3518 <= vdd;
        else
            _3518 <= _3516;
    end
    assign _3733 = _3704[28:28];
    assign _4186 = vdd ? _3733 : _3521;
    assign _4187 = _3739 ? _4186 : _3521;
    assign _4188 = _3745 ? _3521 : _4187;
    assign _4189 = _3751 ? _3521 : _4188;
    assign _4190 = _3755 ? _3521 : _4189;
    assign _4191 = _3759 ? _3521 : _4190;
    assign _4192 = _3775 ? _3521 : _4191;
    assign _4193 = _3790 ? _3521 : _4192;
    assign _4194 = _2608 == _2603;
    assign _4195 = _4194 ? _4193 : _3521;
    assign _3519 = _4195;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3521 <= vdd;
        else
            _3521 <= _3519;
    end
    assign _3734 = _3704[29:29];
    assign _4176 = vdd ? _3734 : _3524;
    assign _4177 = _3739 ? _4176 : _3524;
    assign _4178 = _3745 ? _3524 : _4177;
    assign _4179 = _3751 ? _3524 : _4178;
    assign _4180 = _3755 ? _3524 : _4179;
    assign _4181 = _3759 ? _3524 : _4180;
    assign _4182 = _3775 ? _3524 : _4181;
    assign _4183 = _3790 ? _3524 : _4182;
    assign _4184 = _2608 == _2603;
    assign _4185 = _4184 ? _4183 : _3524;
    assign _3522 = _4185;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3524 <= vdd;
        else
            _3524 <= _3522;
    end
    assign _3735 = _3704[30:30];
    assign _4166 = vdd ? _3735 : _3527;
    assign _4167 = _3739 ? _4166 : _3527;
    assign _4168 = _3745 ? _3527 : _4167;
    assign _4169 = _3751 ? _3527 : _4168;
    assign _4170 = _3755 ? _3527 : _4169;
    assign _4171 = _3759 ? _3527 : _4170;
    assign _4172 = _3775 ? _3527 : _4171;
    assign _4173 = _3790 ? _3527 : _4172;
    assign _4174 = _2608 == _2603;
    assign _4175 = _4174 ? _4173 : _3527;
    assign _3525 = _4175;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3527 <= vdd;
        else
            _3527 <= _3525;
    end
    assign _3736 = _3704[31:31];
    assign _4156 = vdd ? _3736 : _3530;
    assign _4157 = _3739 ? _4156 : _3530;
    assign _4158 = _3745 ? _3530 : _4157;
    assign _4159 = _3751 ? _3530 : _4158;
    assign _4160 = _3755 ? _3530 : _4159;
    assign _4161 = _3759 ? _3530 : _4160;
    assign _4162 = _3775 ? _3530 : _4161;
    assign _4163 = _3790 ? _3530 : _4162;
    assign _4164 = _2608 == _2603;
    assign _4165 = _4164 ? _4163 : _3530;
    assign _3528 = _4165;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3530 <= vdd;
        else
            _3530 <= _3528;
    end
    assign _3531 = { _3530, _3527, _3524, _3521, _3518, _3515, _3512, _3509, _3506, _3503, _3500, _3497, _3494, _3491, _3488, _3485, _3482, _3479, _3476, _3473, _3470, _3467, _3464, _3461, _3458, _3455, _3452, _3449, _3446, _3443, _3440, _3437 };
    assign _3661 = _3434 & _3531;
    assign _4525 = _3667 ? _3661 : _3434;
    assign _4526 = _3671 ? _3434 : _4525;
    assign _4527 = _3357 ? _3434 : _4526;
    assign _4528 = _3349 ? _3434 : _4527;
    assign _3953 = _3538 - _3952;
    assign _3955 = _3953 == _3954;
    assign _4523 = _3955 ? _3951 : _4522;
    assign _3970 = irq[0:0];
    assign _3971 = _38[0:0];
    assign _3972 = _3401[0:0];
    assign _3973 = _3972 & _3971;
    assign _3974 = _3973 | _3970;
    assign _4522 = vdd ? _3974 : gnd;
    assign _3701 = instr[46:46];
    assign _3702 = vdd & vdd;
    assign _3703 = _3702 & _3701;
    assign _4134 = _3703 ? _3685 : _4133;
    assign _4135 = _3739 ? _4133 : _4134;
    assign _4136 = _3745 ? _4133 : _4135;
    assign _4137 = _3751 ? _4133 : _4136;
    assign _4138 = _3755 ? _4133 : _4137;
    assign _4139 = _3759 ? _4133 : _4138;
    assign _4140 = _3775 ? _4133 : _4139;
    assign _4141 = _3790 ? _4133 : _4140;
    assign _3950 = _3538 - _3949;
    assign _4133 = _3960 ? _3950 : _3538;
    assign _4142 = _2608 == _2603;
    assign _4143 = _4142 ? _4141 : _4133;
    assign _3536 = _4143;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3538 <= _3535;
        else
            _3538 <= _3536;
    end
    assign _3957 = _3538 == _3956;
    assign _3958 = ~ _3957;
    assign _3959 = vdd & vdd;
    assign _3960 = _3959 & _3958;
    assign _4524 = _3960 ? _4523 : _4522;
    assign _3402 = _4524;
    assign _3782 = ~ _3397;
    assign _3783 = ~ _3440;
    assign _3784 = vdd & _3783;
    assign _3785 = _3784 & _3782;
    assign _4507 = _3785 ? _3781 : _4506;
    assign _4508 = _3329 ? _4507 : _4506;
    assign _4509 = pcpi_int_ready ? _4506 : _4508;
    assign _4510 = vdd ? _4509 : _4506;
    assign _3777 = ~ _3397;
    assign _3778 = ~ _3440;
    assign _3779 = vdd & _3778;
    assign _3780 = _3779 & _3777;
    assign _4511 = _3780 ? _3776 : _4506;
    assign _4512 = vdd ? _4510 : _4511;
    assign _4513 = _3790 ? _4512 : _4506;
    assign _4531 = _3671 ? _3669 : _3397;
    assign _4532 = _3357 ? _3397 : _4531;
    assign _4533 = _3349 ? _3397 : _4532;
    assign _4534 = _3745 ? _3742 : _3397;
    assign _4535 = _3751 ? _3397 : _4534;
    assign _4536 = _3755 ? _3397 : _4535;
    assign _4537 = _3759 ? _3397 : _4536;
    assign _4538 = _3775 ? _3397 : _4537;
    assign _4539 = _3790 ? _3397 : _4538;
    assign _4540 = _2608 == _2603;
    assign _4541 = _4540 ? _4539 : _3397;
    assign _4542 = _2608 == _2605;
    assign _4543 = _4542 ? _4533 : _4541;
    assign _3395 = _4543;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3397 <= _3394;
        else
            _3397 <= _3395;
    end
    assign _3797 = ~ _3397;
    assign _3241 = _3065[35:35];
    assign _3242 = _2675 & _3241;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3245 <= _3243;
        else
            if (_3242)
                _3245 <= _2674;
    end
    assign _3236 = _3065[34:34];
    assign _3237 = _2675 & _3236;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3240 <= _3238;
        else
            if (_3237)
                _3240 <= _2674;
    end
    assign _3231 = _3065[33:33];
    assign _3232 = _2675 & _3231;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3235 <= _3233;
        else
            if (_3232)
                _3235 <= _2674;
    end
    assign _3226 = _3065[32:32];
    assign _3227 = _2675 & _3226;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3230 <= _3228;
        else
            if (_3227)
                _3230 <= _2674;
    end
    assign _3221 = _3065[31:31];
    assign _3222 = _2675 & _3221;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3225 <= _3223;
        else
            if (_3222)
                _3225 <= _2674;
    end
    assign _3216 = _3065[30:30];
    assign _3217 = _2675 & _3216;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3220 <= _3218;
        else
            if (_3217)
                _3220 <= _2674;
    end
    assign _3211 = _3065[29:29];
    assign _3212 = _2675 & _3211;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3215 <= _3213;
        else
            if (_3212)
                _3215 <= _2674;
    end
    assign _3206 = _3065[28:28];
    assign _3207 = _2675 & _3206;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3210 <= _3208;
        else
            if (_3207)
                _3210 <= _2674;
    end
    assign _3201 = _3065[27:27];
    assign _3202 = _2675 & _3201;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3205 <= _3203;
        else
            if (_3202)
                _3205 <= _2674;
    end
    assign _3196 = _3065[26:26];
    assign _3197 = _2675 & _3196;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3200 <= _3198;
        else
            if (_3197)
                _3200 <= _2674;
    end
    assign _3191 = _3065[25:25];
    assign _3192 = _2675 & _3191;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3195 <= _3193;
        else
            if (_3192)
                _3195 <= _2674;
    end
    assign _3186 = _3065[24:24];
    assign _3187 = _2675 & _3186;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3190 <= _3188;
        else
            if (_3187)
                _3190 <= _2674;
    end
    assign _3181 = _3065[23:23];
    assign _3182 = _2675 & _3181;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3185 <= _3183;
        else
            if (_3182)
                _3185 <= _2674;
    end
    assign _3176 = _3065[22:22];
    assign _3177 = _2675 & _3176;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3180 <= _3178;
        else
            if (_3177)
                _3180 <= _2674;
    end
    assign _3171 = _3065[21:21];
    assign _3172 = _2675 & _3171;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3175 <= _3173;
        else
            if (_3172)
                _3175 <= _2674;
    end
    assign _3166 = _3065[20:20];
    assign _3167 = _2675 & _3166;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3170 <= _3168;
        else
            if (_3167)
                _3170 <= _2674;
    end
    assign _3161 = _3065[19:19];
    assign _3162 = _2675 & _3161;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3165 <= _3163;
        else
            if (_3162)
                _3165 <= _2674;
    end
    assign _3156 = _3065[18:18];
    assign _3157 = _2675 & _3156;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3160 <= _3158;
        else
            if (_3157)
                _3160 <= _2674;
    end
    assign _3151 = _3065[17:17];
    assign _3152 = _2675 & _3151;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3155 <= _3153;
        else
            if (_3152)
                _3155 <= _2674;
    end
    assign _3146 = _3065[16:16];
    assign _3147 = _2675 & _3146;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3150 <= _3148;
        else
            if (_3147)
                _3150 <= _2674;
    end
    assign _3141 = _3065[15:15];
    assign _3142 = _2675 & _3141;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3145 <= _3143;
        else
            if (_3142)
                _3145 <= _2674;
    end
    assign _3136 = _3065[14:14];
    assign _3137 = _2675 & _3136;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3140 <= _3138;
        else
            if (_3137)
                _3140 <= _2674;
    end
    assign _3131 = _3065[13:13];
    assign _3132 = _2675 & _3131;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3135 <= _3133;
        else
            if (_3132)
                _3135 <= _2674;
    end
    assign _3126 = _3065[12:12];
    assign _3127 = _2675 & _3126;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3130 <= _3128;
        else
            if (_3127)
                _3130 <= _2674;
    end
    assign _3121 = _3065[11:11];
    assign _3122 = _2675 & _3121;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3125 <= _3123;
        else
            if (_3122)
                _3125 <= _2674;
    end
    assign _3116 = _3065[10:10];
    assign _3117 = _2675 & _3116;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3120 <= _3118;
        else
            if (_3117)
                _3120 <= _2674;
    end
    assign _3111 = _3065[9:9];
    assign _3112 = _2675 & _3111;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3115 <= _3113;
        else
            if (_3112)
                _3115 <= _2674;
    end
    assign _3106 = _3065[8:8];
    assign _3107 = _2675 & _3106;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3110 <= _3108;
        else
            if (_3107)
                _3110 <= _2674;
    end
    assign _3101 = _3065[7:7];
    assign _3102 = _2675 & _3101;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3105 <= _3103;
        else
            if (_3102)
                _3105 <= _2674;
    end
    assign _3096 = _3065[6:6];
    assign _3097 = _2675 & _3096;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3100 <= _3098;
        else
            if (_3097)
                _3100 <= _2674;
    end
    assign _3091 = _3065[5:5];
    assign _3092 = _2675 & _3091;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3095 <= _3093;
        else
            if (_3092)
                _3095 <= _2674;
    end
    assign _3086 = _3065[4:4];
    assign _3087 = _2675 & _3086;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3090 <= _3088;
        else
            if (_3087)
                _3090 <= _2674;
    end
    assign _3081 = _3065[3:3];
    assign _3082 = _2675 & _3081;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3085 <= _3083;
        else
            if (_3082)
                _3085 <= _2674;
    end
    assign _3076 = _3065[2:2];
    assign _3077 = _2675 & _3076;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3080 <= _3078;
        else
            if (_3077)
                _3080 <= _2674;
    end
    assign _2682 = ~ _2676;
    assign _2685 = _2683 & _2682;
    assign _2693 = _2689 & _2685;
    assign _2713 = _2705 & _2693;
    assign _2761 = _2745 & _2713;
    assign _2873 = _2841 & _2761;
    assign _2683 = ~ _2677;
    assign _2684 = _2683 & _2676;
    assign _2692 = _2689 & _2684;
    assign _2712 = _2705 & _2692;
    assign _2760 = _2745 & _2712;
    assign _2872 = _2841 & _2760;
    assign _2686 = ~ _2676;
    assign _2688 = _2677 & _2686;
    assign _2691 = _2689 & _2688;
    assign _2711 = _2705 & _2691;
    assign _2759 = _2745 & _2711;
    assign _2871 = _2841 & _2759;
    assign _2687 = _2677 & _2676;
    assign _2689 = ~ _2678;
    assign _2690 = _2689 & _2687;
    assign _2710 = _2705 & _2690;
    assign _2758 = _2745 & _2710;
    assign _2870 = _2841 & _2758;
    assign _2694 = ~ _2676;
    assign _2697 = _2695 & _2694;
    assign _2704 = _2678 & _2697;
    assign _2709 = _2705 & _2704;
    assign _2757 = _2745 & _2709;
    assign _2869 = _2841 & _2757;
    assign _2695 = ~ _2677;
    assign _2696 = _2695 & _2676;
    assign _2703 = _2678 & _2696;
    assign _2708 = _2705 & _2703;
    assign _2756 = _2745 & _2708;
    assign _2868 = _2841 & _2756;
    assign _2698 = ~ _2676;
    assign _2700 = _2677 & _2698;
    assign _2702 = _2678 & _2700;
    assign _2707 = _2705 & _2702;
    assign _2755 = _2745 & _2707;
    assign _2867 = _2841 & _2755;
    assign _2699 = _2677 & _2676;
    assign _2701 = _2678 & _2699;
    assign _2705 = ~ _2679;
    assign _2706 = _2705 & _2701;
    assign _2754 = _2745 & _2706;
    assign _2866 = _2841 & _2754;
    assign _2714 = ~ _2676;
    assign _2717 = _2715 & _2714;
    assign _2725 = _2721 & _2717;
    assign _2744 = _2679 & _2725;
    assign _2753 = _2745 & _2744;
    assign _2865 = _2841 & _2753;
    assign _2715 = ~ _2677;
    assign _2716 = _2715 & _2676;
    assign _2724 = _2721 & _2716;
    assign _2743 = _2679 & _2724;
    assign _2752 = _2745 & _2743;
    assign _2864 = _2841 & _2752;
    assign _2718 = ~ _2676;
    assign _2720 = _2677 & _2718;
    assign _2723 = _2721 & _2720;
    assign _2742 = _2679 & _2723;
    assign _2751 = _2745 & _2742;
    assign _2863 = _2841 & _2751;
    assign _2719 = _2677 & _2676;
    assign _2721 = ~ _2678;
    assign _2722 = _2721 & _2719;
    assign _2741 = _2679 & _2722;
    assign _2750 = _2745 & _2741;
    assign _2862 = _2841 & _2750;
    assign _2726 = ~ _2676;
    assign _2729 = _2727 & _2726;
    assign _2736 = _2678 & _2729;
    assign _2740 = _2679 & _2736;
    assign _2749 = _2745 & _2740;
    assign _2861 = _2841 & _2749;
    assign _2727 = ~ _2677;
    assign _2728 = _2727 & _2676;
    assign _2735 = _2678 & _2728;
    assign _2739 = _2679 & _2735;
    assign _2748 = _2745 & _2739;
    assign _2860 = _2841 & _2748;
    assign _2730 = ~ _2676;
    assign _2732 = _2677 & _2730;
    assign _2734 = _2678 & _2732;
    assign _2738 = _2679 & _2734;
    assign _2747 = _2745 & _2738;
    assign _2859 = _2841 & _2747;
    assign _2731 = _2677 & _2676;
    assign _2733 = _2678 & _2731;
    assign _2737 = _2679 & _2733;
    assign _2745 = ~ _2680;
    assign _2746 = _2745 & _2737;
    assign _2858 = _2841 & _2746;
    assign _2762 = ~ _2676;
    assign _2765 = _2763 & _2762;
    assign _2773 = _2769 & _2765;
    assign _2793 = _2785 & _2773;
    assign _2840 = _2680 & _2793;
    assign _2857 = _2841 & _2840;
    assign _2763 = ~ _2677;
    assign _2764 = _2763 & _2676;
    assign _2772 = _2769 & _2764;
    assign _2792 = _2785 & _2772;
    assign _2839 = _2680 & _2792;
    assign _2856 = _2841 & _2839;
    assign _2766 = ~ _2676;
    assign _2768 = _2677 & _2766;
    assign _2771 = _2769 & _2768;
    assign _2791 = _2785 & _2771;
    assign _2838 = _2680 & _2791;
    assign _2855 = _2841 & _2838;
    assign _2767 = _2677 & _2676;
    assign _2769 = ~ _2678;
    assign _2770 = _2769 & _2767;
    assign _2790 = _2785 & _2770;
    assign _2837 = _2680 & _2790;
    assign _2854 = _2841 & _2837;
    assign _2774 = ~ _2676;
    assign _2777 = _2775 & _2774;
    assign _2784 = _2678 & _2777;
    assign _2789 = _2785 & _2784;
    assign _2836 = _2680 & _2789;
    assign _2853 = _2841 & _2836;
    assign _2775 = ~ _2677;
    assign _2776 = _2775 & _2676;
    assign _2783 = _2678 & _2776;
    assign _2788 = _2785 & _2783;
    assign _2835 = _2680 & _2788;
    assign _2852 = _2841 & _2835;
    assign _2778 = ~ _2676;
    assign _2780 = _2677 & _2778;
    assign _2782 = _2678 & _2780;
    assign _2787 = _2785 & _2782;
    assign _2834 = _2680 & _2787;
    assign _2851 = _2841 & _2834;
    assign _2779 = _2677 & _2676;
    assign _2781 = _2678 & _2779;
    assign _2785 = ~ _2679;
    assign _2786 = _2785 & _2781;
    assign _2833 = _2680 & _2786;
    assign _2850 = _2841 & _2833;
    assign _2794 = ~ _2676;
    assign _2797 = _2795 & _2794;
    assign _2805 = _2801 & _2797;
    assign _2824 = _2679 & _2805;
    assign _2832 = _2680 & _2824;
    assign _2849 = _2841 & _2832;
    assign _2795 = ~ _2677;
    assign _2796 = _2795 & _2676;
    assign _2804 = _2801 & _2796;
    assign _2823 = _2679 & _2804;
    assign _2831 = _2680 & _2823;
    assign _2848 = _2841 & _2831;
    assign _2798 = ~ _2676;
    assign _2800 = _2677 & _2798;
    assign _2803 = _2801 & _2800;
    assign _2822 = _2679 & _2803;
    assign _2830 = _2680 & _2822;
    assign _2847 = _2841 & _2830;
    assign _2799 = _2677 & _2676;
    assign _2801 = ~ _2678;
    assign _2802 = _2801 & _2799;
    assign _2821 = _2679 & _2802;
    assign _2829 = _2680 & _2821;
    assign _2846 = _2841 & _2829;
    assign _2806 = ~ _2676;
    assign _2809 = _2807 & _2806;
    assign _2816 = _2678 & _2809;
    assign _2820 = _2679 & _2816;
    assign _2828 = _2680 & _2820;
    assign _2845 = _2841 & _2828;
    assign _2807 = ~ _2677;
    assign _2808 = _2807 & _2676;
    assign _2815 = _2678 & _2808;
    assign _2819 = _2679 & _2815;
    assign _2827 = _2680 & _2819;
    assign _2844 = _2841 & _2827;
    assign _2810 = ~ _2676;
    assign _2812 = _2677 & _2810;
    assign _2814 = _2678 & _2812;
    assign _2818 = _2679 & _2814;
    assign _2826 = _2680 & _2818;
    assign _2843 = _2841 & _2826;
    assign _2811 = _2677 & _2676;
    assign _2813 = _2678 & _2811;
    assign _2817 = _2679 & _2813;
    assign _2825 = _2680 & _2817;
    assign _2841 = ~ _2681;
    assign _2842 = _2841 & _2825;
    assign _2874 = ~ _2676;
    assign _2877 = _2875 & _2874;
    assign _2885 = _2881 & _2877;
    assign _2905 = _2897 & _2885;
    assign _2953 = _2937 & _2905;
    assign _3064 = _2681 & _2953;
    assign _2875 = ~ _2677;
    assign _2876 = _2875 & _2676;
    assign _2884 = _2881 & _2876;
    assign _2904 = _2897 & _2884;
    assign _2952 = _2937 & _2904;
    assign _3063 = _2681 & _2952;
    assign _2878 = ~ _2676;
    assign _2880 = _2677 & _2878;
    assign _2883 = _2881 & _2880;
    assign _2903 = _2897 & _2883;
    assign _2951 = _2937 & _2903;
    assign _3062 = _2681 & _2951;
    assign _2879 = _2677 & _2676;
    assign _2881 = ~ _2678;
    assign _2882 = _2881 & _2879;
    assign _2902 = _2897 & _2882;
    assign _2950 = _2937 & _2902;
    assign _3061 = _2681 & _2950;
    assign _2886 = ~ _2676;
    assign _2889 = _2887 & _2886;
    assign _2896 = _2678 & _2889;
    assign _2901 = _2897 & _2896;
    assign _2949 = _2937 & _2901;
    assign _3060 = _2681 & _2949;
    assign _2887 = ~ _2677;
    assign _2888 = _2887 & _2676;
    assign _2895 = _2678 & _2888;
    assign _2900 = _2897 & _2895;
    assign _2948 = _2937 & _2900;
    assign _3059 = _2681 & _2948;
    assign _2890 = ~ _2676;
    assign _2892 = _2677 & _2890;
    assign _2894 = _2678 & _2892;
    assign _2899 = _2897 & _2894;
    assign _2947 = _2937 & _2899;
    assign _3058 = _2681 & _2947;
    assign _2891 = _2677 & _2676;
    assign _2893 = _2678 & _2891;
    assign _2897 = ~ _2679;
    assign _2898 = _2897 & _2893;
    assign _2946 = _2937 & _2898;
    assign _3057 = _2681 & _2946;
    assign _2906 = ~ _2676;
    assign _2909 = _2907 & _2906;
    assign _2917 = _2913 & _2909;
    assign _2936 = _2679 & _2917;
    assign _2945 = _2937 & _2936;
    assign _3056 = _2681 & _2945;
    assign _2907 = ~ _2677;
    assign _2908 = _2907 & _2676;
    assign _2916 = _2913 & _2908;
    assign _2935 = _2679 & _2916;
    assign _2944 = _2937 & _2935;
    assign _3055 = _2681 & _2944;
    assign _2910 = ~ _2676;
    assign _2912 = _2677 & _2910;
    assign _2915 = _2913 & _2912;
    assign _2934 = _2679 & _2915;
    assign _2943 = _2937 & _2934;
    assign _3054 = _2681 & _2943;
    assign _2911 = _2677 & _2676;
    assign _2913 = ~ _2678;
    assign _2914 = _2913 & _2911;
    assign _2933 = _2679 & _2914;
    assign _2942 = _2937 & _2933;
    assign _3053 = _2681 & _2942;
    assign _2918 = ~ _2676;
    assign _2921 = _2919 & _2918;
    assign _2928 = _2678 & _2921;
    assign _2932 = _2679 & _2928;
    assign _2941 = _2937 & _2932;
    assign _3052 = _2681 & _2941;
    assign _2919 = ~ _2677;
    assign _2920 = _2919 & _2676;
    assign _2927 = _2678 & _2920;
    assign _2931 = _2679 & _2927;
    assign _2940 = _2937 & _2931;
    assign _3051 = _2681 & _2940;
    assign _2922 = ~ _2676;
    assign _2924 = _2677 & _2922;
    assign _2926 = _2678 & _2924;
    assign _2930 = _2679 & _2926;
    assign _2939 = _2937 & _2930;
    assign _3050 = _2681 & _2939;
    assign _2923 = _2677 & _2676;
    assign _2925 = _2678 & _2923;
    assign _2929 = _2679 & _2925;
    assign _2937 = ~ _2680;
    assign _2938 = _2937 & _2929;
    assign _3049 = _2681 & _2938;
    assign _2954 = ~ _2676;
    assign _2957 = _2955 & _2954;
    assign _2965 = _2961 & _2957;
    assign _2985 = _2977 & _2965;
    assign _3032 = _2680 & _2985;
    assign _3048 = _2681 & _3032;
    assign _2955 = ~ _2677;
    assign _2956 = _2955 & _2676;
    assign _2964 = _2961 & _2956;
    assign _2984 = _2977 & _2964;
    assign _3031 = _2680 & _2984;
    assign _3047 = _2681 & _3031;
    assign _2958 = ~ _2676;
    assign _2960 = _2677 & _2958;
    assign _2963 = _2961 & _2960;
    assign _2983 = _2977 & _2963;
    assign _3030 = _2680 & _2983;
    assign _3046 = _2681 & _3030;
    assign _2959 = _2677 & _2676;
    assign _2961 = ~ _2678;
    assign _2962 = _2961 & _2959;
    assign _2982 = _2977 & _2962;
    assign _3029 = _2680 & _2982;
    assign _3045 = _2681 & _3029;
    assign _2966 = ~ _2676;
    assign _2969 = _2967 & _2966;
    assign _2976 = _2678 & _2969;
    assign _2981 = _2977 & _2976;
    assign _3028 = _2680 & _2981;
    assign _3044 = _2681 & _3028;
    assign _2967 = ~ _2677;
    assign _2968 = _2967 & _2676;
    assign _2975 = _2678 & _2968;
    assign _2980 = _2977 & _2975;
    assign _3027 = _2680 & _2980;
    assign _3043 = _2681 & _3027;
    assign _2970 = ~ _2676;
    assign _2972 = _2677 & _2970;
    assign _2974 = _2678 & _2972;
    assign _2979 = _2977 & _2974;
    assign _3026 = _2680 & _2979;
    assign _3042 = _2681 & _3026;
    assign _2971 = _2677 & _2676;
    assign _2973 = _2678 & _2971;
    assign _2977 = ~ _2679;
    assign _2978 = _2977 & _2973;
    assign _3025 = _2680 & _2978;
    assign _3041 = _2681 & _3025;
    assign _2986 = ~ _2676;
    assign _2989 = _2987 & _2986;
    assign _2997 = _2993 & _2989;
    assign _3016 = _2679 & _2997;
    assign _3024 = _2680 & _3016;
    assign _3040 = _2681 & _3024;
    assign _2987 = ~ _2677;
    assign _2988 = _2987 & _2676;
    assign _2996 = _2993 & _2988;
    assign _3015 = _2679 & _2996;
    assign _3023 = _2680 & _3015;
    assign _3039 = _2681 & _3023;
    assign _2990 = ~ _2676;
    assign _2992 = _2677 & _2990;
    assign _2995 = _2993 & _2992;
    assign _3014 = _2679 & _2995;
    assign _3022 = _2680 & _3014;
    assign _3038 = _2681 & _3022;
    assign _2991 = _2677 & _2676;
    assign _2993 = ~ _2678;
    assign _2994 = _2993 & _2991;
    assign _3013 = _2679 & _2994;
    assign _3021 = _2680 & _3013;
    assign _3037 = _2681 & _3021;
    assign _2998 = ~ _2676;
    assign _3001 = _2999 & _2998;
    assign _3008 = _2678 & _3001;
    assign _3012 = _2679 & _3008;
    assign _3020 = _2680 & _3012;
    assign _3036 = _2681 & _3020;
    assign _2999 = ~ _2677;
    assign _3000 = _2999 & _2676;
    assign _3007 = _2678 & _3000;
    assign _3011 = _2679 & _3007;
    assign _3019 = _2680 & _3011;
    assign _3035 = _2681 & _3019;
    assign _3002 = ~ _2676;
    assign _3004 = _2677 & _3002;
    assign _3006 = _2678 & _3004;
    assign _3010 = _2679 & _3006;
    assign _3018 = _2680 & _3010;
    assign _3034 = _2681 & _3018;
    assign _2676 = _2672[0:0];
    assign _2677 = _2672[1:1];
    assign _3003 = _2677 & _2676;
    assign _2678 = _2672[2:2];
    assign _3005 = _2678 & _3003;
    assign _2679 = _2672[3:3];
    assign _3009 = _2679 & _3005;
    assign _2680 = _2672[4:4];
    assign _3017 = _2680 & _3009;
    assign _3565 = _3393[0:0];
    assign _3570 = { _3568, _3565 };
    assign _3572 = _3571 | _3570;
    assign _3564 = _3393[0:0];
    assign _4978 = _3564 ? _3563 : _3562;
    assign _4979 = vdd ? _3572 : _4978;
    assign _4980 = _3654 ? _4979 : decoded_rd;
    assign _3748 = _2672 | _3747;
    assign _4981 = _3751 ? _3748 : _2672;
    assign _4982 = _3755 ? _2672 : _4981;
    assign _4983 = _3759 ? _2672 : _4982;
    assign _4984 = _3775 ? _2672 : _4983;
    assign _4985 = _3790 ? _2672 : _4984;
    assign _4986 = _3813 ? _3812 : _2672;
    assign _4987 = _2608 == _2601;
    assign _4988 = _4987 ? _4986 : _2672;
    assign _4989 = _2608 == _2603;
    assign _4990 = _4989 ? _4985 : _4988;
    assign _4991 = _2608 == _2605;
    assign _4992 = _4991 ? _4980 : _4990;
    assign _2670 = _4992;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2672 <= _2669;
        else
            _2672 <= _2670;
    end
    assign _2681 = _2672[5:5];
    assign _3033 = _2681 & _3017;
    assign _3065 = { _3033, _3034, _3035, _3036, _3037, _3038, _3039, _3040, _3041, _3042, _3043, _3044, _3045, _3046, _3047, _3048, _3049, _3050, _3051, _3052, _3053, _3054, _3055, _3056, _3057, _3058, _3059, _3060, _3061, _3062, _3063, _3064, _2842, _2843, _2844, _2845, _2846, _2847, _2848, _2849, _2850, _2851, _2852, _2853, _2854, _2855, _2856, _2857, _2858, _2859, _2860, _2861, _2862, _2863, _2864, _2865, _2866, _2867, _2868, _2869, _2870, _2871, _2872, _2873 };
    assign _3071 = _3065[1:1];
    assign _4958 = vdd ? vdd : gnd;
    assign _4959 = vdd ? vdd : gnd;
    assign _4960 = vdd ? vdd : gnd;
    assign _4961 = vdd ? vdd : gnd;
    assign _3666 = _3393[1:1];
    assign _3667 = vdd & _3666;
    assign _4962 = _3667 ? _4961 : gnd;
    assign _3576 = _3393 == _3575;
    assign _3577 = _3576 ? _3574 : _3573;
    assign _3580 = _3393 == _3579;
    assign _3581 = _3580 ? _3578 : _3577;
    assign _4544 = _3654 ? _3581 : _3393;
    assign _4545 = _2608 == _2605;
    assign _4546 = _4545 ? _4544 : _3393;
    assign _3391 = _4546;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3393 <= _3390;
        else
            _3393 <= _3391;
    end
    assign _3670 = _3393[0:0];
    assign _3671 = vdd & _3670;
    assign _4963 = _3671 ? _4960 : _4962;
    assign _4964 = _3357 ? _4959 : _4963;
    assign _4965 = _3349 ? _4958 : _4964;
    assign _4966 = _2608 == _2605;
    assign _4967 = _4966 ? _4965 : gnd;
    assign _2675 = _4967;
    assign _3072 = _2675 & _3071;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3075 <= _3073;
        else
            if (_3072)
                _3075 <= _2674;
    end
    always @* begin
        case (decoded_rs1)
        0: _3247 <= _3070;
        1: _3247 <= _3075;
        2: _3247 <= _3080;
        3: _3247 <= _3085;
        4: _3247 <= _3090;
        5: _3247 <= _3095;
        6: _3247 <= _3100;
        7: _3247 <= _3105;
        8: _3247 <= _3110;
        9: _3247 <= _3115;
        10: _3247 <= _3120;
        11: _3247 <= _3125;
        12: _3247 <= _3130;
        13: _3247 <= _3135;
        14: _3247 <= _3140;
        15: _3247 <= _3145;
        16: _3247 <= _3150;
        17: _3247 <= _3155;
        18: _3247 <= _3160;
        19: _3247 <= _3165;
        20: _3247 <= _3170;
        21: _3247 <= _3175;
        22: _3247 <= _3180;
        23: _3247 <= _3185;
        24: _3247 <= _3190;
        25: _3247 <= _3195;
        26: _3247 <= _3200;
        27: _3247 <= _3205;
        28: _3247 <= _3210;
        29: _3247 <= _3215;
        30: _3247 <= _3220;
        31: _3247 <= _3225;
        32: _3247 <= _3230;
        33: _3247 <= _3235;
        34: _3247 <= _3240;
        default: _3247 <= _3245;
        endcase
    end
    assign _3683 = decoded_rs1 == _3682;
    assign _3684 = ~ _3683;
    assign _3685 = _3684 ? _3247 : _3681;
    assign _3704 = _3685 | _37;
    assign _3706 = _3704[1:1];
    assign _4456 = vdd ? _3706 : _3440;
    assign _3738 = instr[44:44];
    assign _3739 = vdd & _3738;
    assign _4457 = _3739 ? _4456 : _3440;
    assign _4458 = _3745 ? _3440 : _4457;
    assign _4459 = _3751 ? _3440 : _4458;
    assign _4460 = _3755 ? _3440 : _4459;
    assign _4461 = _3759 ? _3440 : _4460;
    assign _4462 = _3775 ? _3440 : _4461;
    assign _4463 = _3790 ? _3440 : _4462;
    assign _4464 = _2608 == _2603;
    assign _4465 = _4464 ? _4463 : _3440;
    assign _3438 = _4465;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3440 <= vdd;
        else
            _3440 <= _3438;
    end
    assign _3798 = ~ _3440;
    assign _3799 = vdd & _3798;
    assign _3800 = _3799 & _3797;
    assign _4514 = _3800 ? _3796 : _4506;
    assign _3967 = _3333 - _3966;
    assign _4947 = _3333[0:0];
    assign _4948 = _3333[1:1];
    assign _4949 = _3333[2:2];
    assign _4950 = _3333[3:3];
    assign _4951 = _4950 | _4949;
    assign _4952 = _4951 | _4948;
    assign _4953 = _4952 | _4947;
    assign _4954 = _4953 ? _3967 : _3333;
    assign _3968 = ~ pcpi_int_wait;
    assign _5160 = pcpi_int_ready ? _3786 : _3789;
    assign _5161 = vdd ? _5160 : _2632;
    assign _5162 = vdd ? _5161 : _2632;
    assign _5163 = _3790 ? _5162 : _2632;
    assign _5164 = pcpi_int_ready ? _3801 : _3803;
    assign _5165 = _3805 ? _5164 : _2632;
    assign _5166 = _2608 == _2602;
    assign _5167 = _5166 ? _5165 : _2632;
    assign _5168 = _2608 == _2603;
    assign _5169 = _5168 ? _5163 : _5167;
    assign _2630 = _5169;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2632 <= _2629;
        else
            _2632 <= _2630;
    end
    assign _3969 = _2632 & _3968;
    assign _4955 = _3969 ? _4954 : _3965;
    assign _4956 = vdd ? _4955 : _3333;
    assign _3331 = _4956;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3333 <= _3330;
        else
            _3333 <= _3331;
    end
    assign _3964 = _3333 == _3963;
    assign _4957 = vdd ? _3964 : _3329;
    assign _3327 = _4957;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3329 <= _3326;
        else
            _3329 <= _3327;
    end
    assign _4515 = _3329 ? _4514 : _4506;
    assign _4516 = pcpi_int_ready ? _4506 : _4515;
    assign _3804 = instr[47:47];
    assign _3805 = vdd & _3804;
    assign _4517 = _3805 ? _4516 : _4506;
    assign _3975 = irq[1:1];
    assign _3976 = _38[1:1];
    assign _3977 = _3401[1:1];
    assign _3978 = _3977 & _3976;
    assign _3979 = _3978 | _3975;
    assign _4506 = vdd ? _3979 : gnd;
    assign _4518 = _2608 == _2602;
    assign _4519 = _4518 ? _4517 : _4506;
    assign _4520 = _2608 == _2603;
    assign _4521 = _4520 ? _4513 : _4519;
    assign _3403 = _4521;
    assign _3980 = irq[2:2];
    assign _3981 = _38[2:2];
    assign _3982 = _3401[2:2];
    assign _3983 = _3982 & _3981;
    assign _3984 = _3983 | _3980;
    assign _4505 = vdd ? _3984 : gnd;
    assign _3404 = _4505;
    assign _3985 = irq[3:3];
    assign _3986 = _38[3:3];
    assign _3987 = _3401[3:3];
    assign _3988 = _3987 & _3986;
    assign _3989 = _3988 | _3985;
    assign _4504 = vdd ? _3989 : gnd;
    assign _3405 = _4504;
    assign _3990 = irq[4:4];
    assign _3991 = _38[4:4];
    assign _3992 = _3401[4:4];
    assign _3993 = _3992 & _3991;
    assign _3994 = _3993 | _3990;
    assign _4503 = vdd ? _3994 : gnd;
    assign _3406 = _4503;
    assign _3995 = irq[5:5];
    assign _3996 = _38[5:5];
    assign _3997 = _3401[5:5];
    assign _3998 = _3997 & _3996;
    assign _3999 = _3998 | _3995;
    assign _4502 = vdd ? _3999 : gnd;
    assign _3407 = _4502;
    assign _4000 = irq[6:6];
    assign _4001 = _38[6:6];
    assign _4002 = _3401[6:6];
    assign _4003 = _4002 & _4001;
    assign _4004 = _4003 | _4000;
    assign _4501 = vdd ? _4004 : gnd;
    assign _3408 = _4501;
    assign _4005 = irq[7:7];
    assign _4006 = _38[7:7];
    assign _4007 = _3401[7:7];
    assign _4008 = _4007 & _4006;
    assign _4009 = _4008 | _4005;
    assign _4500 = vdd ? _4009 : gnd;
    assign _3409 = _4500;
    assign _4010 = irq[8:8];
    assign _4011 = _38[8:8];
    assign _4012 = _3401[8:8];
    assign _4013 = _4012 & _4011;
    assign _4014 = _4013 | _4010;
    assign _4499 = vdd ? _4014 : gnd;
    assign _3410 = _4499;
    assign _4015 = irq[9:9];
    assign _4016 = _38[9:9];
    assign _4017 = _3401[9:9];
    assign _4018 = _4017 & _4016;
    assign _4019 = _4018 | _4015;
    assign _4498 = vdd ? _4019 : gnd;
    assign _3411 = _4498;
    assign _4020 = irq[10:10];
    assign _4021 = _38[10:10];
    assign _4022 = _3401[10:10];
    assign _4023 = _4022 & _4021;
    assign _4024 = _4023 | _4020;
    assign _4497 = vdd ? _4024 : gnd;
    assign _3412 = _4497;
    assign _4025 = irq[11:11];
    assign _4026 = _38[11:11];
    assign _4027 = _3401[11:11];
    assign _4028 = _4027 & _4026;
    assign _4029 = _4028 | _4025;
    assign _4496 = vdd ? _4029 : gnd;
    assign _3413 = _4496;
    assign _4030 = irq[12:12];
    assign _4031 = _38[12:12];
    assign _4032 = _3401[12:12];
    assign _4033 = _4032 & _4031;
    assign _4034 = _4033 | _4030;
    assign _4495 = vdd ? _4034 : gnd;
    assign _3414 = _4495;
    assign _4035 = irq[13:13];
    assign _4036 = _38[13:13];
    assign _4037 = _3401[13:13];
    assign _4038 = _4037 & _4036;
    assign _4039 = _4038 | _4035;
    assign _4494 = vdd ? _4039 : gnd;
    assign _3415 = _4494;
    assign _4040 = irq[14:14];
    assign _4041 = _38[14:14];
    assign _4042 = _3401[14:14];
    assign _4043 = _4042 & _4041;
    assign _4044 = _4043 | _4040;
    assign _4493 = vdd ? _4044 : gnd;
    assign _3416 = _4493;
    assign _4045 = irq[15:15];
    assign _4046 = _38[15:15];
    assign _4047 = _3401[15:15];
    assign _4048 = _4047 & _4046;
    assign _4049 = _4048 | _4045;
    assign _4492 = vdd ? _4049 : gnd;
    assign _3417 = _4492;
    assign _4050 = irq[16:16];
    assign _4051 = _38[16:16];
    assign _4052 = _3401[16:16];
    assign _4053 = _4052 & _4051;
    assign _4054 = _4053 | _4050;
    assign _4491 = vdd ? _4054 : gnd;
    assign _3418 = _4491;
    assign _4055 = irq[17:17];
    assign _4056 = _38[17:17];
    assign _4057 = _3401[17:17];
    assign _4058 = _4057 & _4056;
    assign _4059 = _4058 | _4055;
    assign _4490 = vdd ? _4059 : gnd;
    assign _3419 = _4490;
    assign _4060 = irq[18:18];
    assign _4061 = _38[18:18];
    assign _4062 = _3401[18:18];
    assign _4063 = _4062 & _4061;
    assign _4064 = _4063 | _4060;
    assign _4489 = vdd ? _4064 : gnd;
    assign _3420 = _4489;
    assign _4065 = irq[19:19];
    assign _4066 = _38[19:19];
    assign _4067 = _3401[19:19];
    assign _4068 = _4067 & _4066;
    assign _4069 = _4068 | _4065;
    assign _4488 = vdd ? _4069 : gnd;
    assign _3421 = _4488;
    assign _4070 = irq[20:20];
    assign _4071 = _38[20:20];
    assign _4072 = _3401[20:20];
    assign _4073 = _4072 & _4071;
    assign _4074 = _4073 | _4070;
    assign _4487 = vdd ? _4074 : gnd;
    assign _3422 = _4487;
    assign _4075 = irq[21:21];
    assign _4076 = _38[21:21];
    assign _4077 = _3401[21:21];
    assign _4078 = _4077 & _4076;
    assign _4079 = _4078 | _4075;
    assign _4486 = vdd ? _4079 : gnd;
    assign _3423 = _4486;
    assign _4080 = irq[22:22];
    assign _4081 = _38[22:22];
    assign _4082 = _3401[22:22];
    assign _4083 = _4082 & _4081;
    assign _4084 = _4083 | _4080;
    assign _4485 = vdd ? _4084 : gnd;
    assign _3424 = _4485;
    assign _4085 = irq[23:23];
    assign _4086 = _38[23:23];
    assign _4087 = _3401[23:23];
    assign _4088 = _4087 & _4086;
    assign _4089 = _4088 | _4085;
    assign _4484 = vdd ? _4089 : gnd;
    assign _3425 = _4484;
    assign _4090 = irq[24:24];
    assign _4091 = _38[24:24];
    assign _4092 = _3401[24:24];
    assign _4093 = _4092 & _4091;
    assign _4094 = _4093 | _4090;
    assign _4483 = vdd ? _4094 : gnd;
    assign _3426 = _4483;
    assign _4095 = irq[25:25];
    assign _4096 = _38[25:25];
    assign _4097 = _3401[25:25];
    assign _4098 = _4097 & _4096;
    assign _4099 = _4098 | _4095;
    assign _4482 = vdd ? _4099 : gnd;
    assign _3427 = _4482;
    assign _4100 = irq[26:26];
    assign _4101 = _38[26:26];
    assign _4102 = _3401[26:26];
    assign _4103 = _4102 & _4101;
    assign _4104 = _4103 | _4100;
    assign _4481 = vdd ? _4104 : gnd;
    assign _3428 = _4481;
    assign _4105 = irq[27:27];
    assign _4106 = _38[27:27];
    assign _4107 = _3401[27:27];
    assign _4108 = _4107 & _4106;
    assign _4109 = _4108 | _4105;
    assign _4480 = vdd ? _4109 : gnd;
    assign _3429 = _4480;
    assign _4110 = irq[28:28];
    assign _4111 = _38[28:28];
    assign _4112 = _3401[28:28];
    assign _4113 = _4112 & _4111;
    assign _4114 = _4113 | _4110;
    assign _4479 = vdd ? _4114 : gnd;
    assign _3430 = _4479;
    assign _4115 = irq[29:29];
    assign _4116 = _38[29:29];
    assign _4117 = _3401[29:29];
    assign _4118 = _4117 & _4116;
    assign _4119 = _4118 | _4115;
    assign _4478 = vdd ? _4119 : gnd;
    assign _3431 = _4478;
    assign _4120 = irq[30:30];
    assign _4121 = _38[30:30];
    assign _4122 = _3401[30:30];
    assign _4123 = _4122 & _4121;
    assign _4124 = _4123 | _4120;
    assign _4477 = vdd ? _4124 : gnd;
    assign _3432 = _4477;
    assign _4125 = irq[31:31];
    assign _4126 = _38[31:31];
    assign _4127 = _3401[31:31];
    assign _4128 = _4127 & _4126;
    assign _4129 = _4128 | _4125;
    assign _4476 = vdd ? _4129 : gnd;
    assign _3433 = _4476;
    assign _3434 = { _3433, _3432, _3431, _3430, _3429, _3428, _3427, _3426, _3425, _3424, _3423, _3422, _3421, _3420, _3419, _3418, _3417, _3416, _3415, _3414, _3413, _3412, _3411, _3410, _3409, _3408, _3407, _3406, _3405, _3404, _3403, _3402 };
    assign _4529 = _2608 == _2605;
    assign _4530 = _4529 ? _4528 : _3434;
    assign _3399 = _4530;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3401 <= _3398;
        else
            _3401 <= _3399;
    end
    assign _4910 = _3401[31:31];
    assign _4911 = _4910 | _4909;
    assign _4912 = _4911 | _4908;
    assign _4913 = _4912 | _4907;
    assign _4914 = _4913 | _4906;
    assign _4915 = _4914 | _4905;
    assign _4916 = _4915 | _4904;
    assign _4917 = _4916 | _4903;
    assign _4918 = _4917 | _4902;
    assign _4919 = _4918 | _4901;
    assign _4920 = _4919 | _4900;
    assign _4921 = _4920 | _4899;
    assign _4922 = _4921 | _4898;
    assign _4923 = _4922 | _4897;
    assign _4924 = _4923 | _4896;
    assign _4925 = _4924 | _4895;
    assign _4926 = _4925 | _4894;
    assign _4927 = _4926 | _4893;
    assign _4928 = _4927 | _4892;
    assign _4929 = _4928 | _4891;
    assign _4930 = _4929 | _4890;
    assign _4931 = _4930 | _4889;
    assign _4932 = _4931 | _4888;
    assign _4933 = _4932 | _4887;
    assign _4934 = _4933 | _4886;
    assign _4935 = _4934 | _4885;
    assign _4936 = _4935 | _4884;
    assign _4937 = _4936 | _4883;
    assign _4938 = _4937 | _4882;
    assign _4939 = _4938 | _4881;
    assign _4940 = _4939 | _4880;
    assign _4941 = _4940 | _4879;
    assign _4942 = _4941 ? _3946 : _3553;
    assign _4943 = _3561 ? _4942 : _3946;
    assign _4944 = _3654 ? _3946 : _4943;
    assign _4945 = _2608 == _2605;
    assign _4946 = _4945 ? _4944 : _3946;
    assign _3335 = _4946;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3337 <= _3334;
        else
            _3337 <= _3335;
    end
    assign _3559 = _2628 | _3337;
    assign _3560 = vdd & _3559;
    assign _3561 = _3560 & _3558;
    assign _4857 = _3561 ? _3658 : _4856;
    assign _4858 = _3654 ? _3658 : _4857;
    assign _3744 = instr[43:43];
    assign _3745 = vdd & _3744;
    assign _4859 = _3745 ? _3741 : _3349;
    assign _3749 = instr[42:42];
    assign _3750 = vdd & vdd;
    assign _3751 = _3750 & _3749;
    assign _4860 = _3751 ? _3349 : _4859;
    assign _3753 = instr[41:41];
    assign _3754 = vdd & vdd;
    assign _3755 = _3754 & _3753;
    assign _4861 = _3755 ? _3349 : _4860;
    assign _3759 = is[0:0];
    assign _4862 = _3759 ? _3349 : _4861;
    assign _3775 = is[14:14];
    assign _4863 = _3775 ? _3349 : _4862;
    assign _3790 = instr[47:47];
    assign _4864 = _3790 ? _3349 : _4863;
    assign _3809 = instr[3:3];
    assign _4865 = _3813 ? _3287 : _3809;
    assign _4866 = _2608 == _2601;
    assign _4867 = _4866 ? _4865 : _3349;
    assign _4868 = _2608 == _2603;
    assign _4869 = _4868 ? _4864 : _4867;
    assign _4870 = _2608 == _2605;
    assign _4871 = _4870 ? _4858 : _4869;
    assign _3347 = _4871;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3349 <= _3346;
        else
            _3349 <= _3347;
    end
    assign _4975 = _3349 ? _4968 : _4974;
    assign _4976 = _2608 == _2605;
    assign _4977 = _4976 ? _4975 : _2673;
    assign _2674 = _4977;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3070 <= _3068;
        else
            if (_3067)
                _3070 <= _2674;
    end
    always @* begin
        case (decoded_rs2)
        0: _3246 <= _3070;
        1: _3246 <= _3075;
        2: _3246 <= _3080;
        3: _3246 <= _3085;
        4: _3246 <= _3090;
        5: _3246 <= _3095;
        6: _3246 <= _3100;
        7: _3246 <= _3105;
        8: _3246 <= _3110;
        9: _3246 <= _3115;
        10: _3246 <= _3120;
        11: _3246 <= _3125;
        12: _3246 <= _3130;
        13: _3246 <= _3135;
        14: _3246 <= _3140;
        15: _3246 <= _3145;
        16: _3246 <= _3150;
        17: _3246 <= _3155;
        18: _3246 <= _3160;
        19: _3246 <= _3165;
        20: _3246 <= _3170;
        21: _3246 <= _3175;
        22: _3246 <= _3180;
        23: _3246 <= _3185;
        24: _3246 <= _3190;
        25: _3246 <= _3195;
        26: _3246 <= _3200;
        27: _3246 <= _3205;
        28: _3246 <= _3210;
        29: _3246 <= _3215;
        30: _3246 <= _3220;
        31: _3246 <= _3225;
        32: _3246 <= _3230;
        33: _3246 <= _3235;
        34: _3246 <= _3240;
        default: _3246 <= _3245;
        endcase
    end
    assign _3688 = decoded_rs2 == _3687;
    assign _3689 = ~ _3688;
    assign _3690 = _3689 ? _3246 : _3686;
    assign _3806 = _3690[4:0];
    assign _3840 = _3389 - _3839;
    assign _3816 = _3389 - _3815;
    assign _3867 = _3389 < _3866;
    assign _3868 = ~ _3867;
    assign _4561 = _3868 ? _3840 : _3816;
    assign _4562 = _3870 ? _4131 : _4561;
    assign _4563 = _2608 == _2600;
    assign _4564 = _4563 ? _4562 : _4131;
    assign _4565 = _2608 == _2602;
    assign _4566 = _4565 ? _3806 : _4564;
    assign _4567 = _2608 == _2603;
    assign _4568 = _4567 ? _4560 : _4566;
    assign _3387 = _4568;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3389 <= _3386;
        else
            _3389 <= _3387;
    end
    assign _3870 = _3389 == _3869;
    assign _5003 = _3870 ? _2664 : _5002;
    assign _3877 = _2664 + decoded_imm;
    assign _5139 = mem_done ? _3942 : _2648;
    assign _4152 = _3888 ? _3876 : gnd;
    assign _4153 = _3890 ? _4152 : gnd;
    assign _4154 = _2608 == _2599;
    assign _4155 = _4154 ? _4153 : gnd;
    assign _3532 = _4155;
    assign _5140 = _3532 ? _3939 : _5139;
    assign _2646 = _5140;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2648 <= _2645;
        else
            _2648 <= _2646;
    end
    assign _3888 = ~ _2648;
    assign _5004 = _3888 ? _3877 : _2664;
    assign _3889 = ~ _2636;
    assign _3890 = _3889 | mem_done;
    assign _5005 = _3890 ? _5004 : _2664;
    assign _3917 = _2664 + decoded_imm;
    assign _5141 = mem_done ? _3943 : _2644;
    assign _4148 = _3935 ? _3916 : gnd;
    assign _4149 = _3937 ? _4148 : gnd;
    assign _4150 = _2608 == _2598;
    assign _4151 = _4150 ? _4149 : gnd;
    assign _3533 = _4151;
    assign _5142 = _3533 ? _3940 : _5141;
    assign _2642 = _5142;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2644 <= _2641;
        else
            _2644 <= _2642;
    end
    assign _3935 = ~ _2644;
    assign _5006 = _3935 ? _3917 : _2664;
    assign _5007 = _3937 ? _5006 : _2664;
    assign _5008 = _2608 == _2598;
    assign _5009 = _5008 ? _5007 : _2664;
    assign _5010 = _2608 == _2599;
    assign _5011 = _5010 ? _5005 : _5009;
    assign _5012 = _2608 == _2600;
    assign _5013 = _5012 ? _5003 : _5011;
    assign _5014 = _2608 == _2603;
    assign _5015 = _5014 ? _5001 : _5013;
    assign _2662 = _5015;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2664 <= _2661;
        else
            _2664 <= _2662;
    end
    assign _3248 = _2664 < _2660;
    assign _3259 = is[7:7];
    assign _3279 = _3259 ? _3258 : _3248;
    assign _3262 = instr[9:9];
    assign _3273 = instr[7:7];
    assign _3282 = _3273 | _3262;
    assign _3276 = instr[5:5];
    assign _3278 = instr[4:4];
    assign _3284 = _3278 | _3276;
    assign _3286 = _3284 | _3282;
    assign _3287 = _3286 ? _3285 : _3279;
    assign _4144 = _3287 ? _3810 : gnd;
    assign _3813 = is[9:9];
    assign _4145 = _3813 ? _4144 : gnd;
    assign _4146 = _2608 == _2601;
    assign _4147 = _4146 ? _4145 : gnd;
    assign _3534 = _4147;
    assign _5138 = _3534 ? _3941 : _5137;
    assign _2650 = _5138;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2652 <= _2649;
        else
            _2652 <= _2650;
    end
    assign _3948 = _2652 & mem_done;
    assign _5176 = _2608 == _2598;
    assign _5177 = _5176 ? _5175 : _3948;
    assign _5178 = _2608 == _2599;
    assign _5179 = _5178 ? _5173 : _5177;
    assign _5180 = _2608 == _2601;
    assign _5181 = _5180 ? _5171 : _5179;
    assign _2626 = _5181;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2628 <= _2625;
        else
            _2628 <= _2626;
    end
    assign _3651 = _2628 & _3650;
    assign _3652 = _3651 & _3649;
    assign _3653 = _3652 | _3584;
    assign _3654 = vdd & _3653;
    assign _5156 = _3654 ? _2636 : _5155;
    assign _5157 = _2608 == _2605;
    assign _5158 = _5157 ? _5156 : _2636;
    assign _5159 = mem_done ? _3945 : _5158;
    assign _2634 = _5159;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2636 <= _2633;
        else
            _2636 <= _2634;
    end
    assign _3936 = ~ _2636;
    assign _3937 = _3936 | mem_done;
    assign _5240 = _3937 ? _5239 : _2608;
    assign _5241 = _2608 == _2598;
    assign _5242 = _5241 ? _5240 : _2608;
    assign _5243 = _2608 == _2599;
    assign _5244 = _5243 ? _5238 : _5242;
    assign _5245 = _2608 == _2600;
    assign _5246 = _5245 ? _5236 : _5244;
    assign _5247 = _2608 == _2601;
    assign _5248 = _5247 ? _5235 : _5246;
    assign _5249 = _2608 == _2602;
    assign _5250 = _5249 ? _5233 : _5248;
    assign _5251 = _2608 == _2603;
    assign _5252 = _5251 ? _5227 : _5250;
    assign _5253 = _2608 == _2605;
    assign _5254 = _5253 ? _5207 : _5252;
    assign _2606 = _5254;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2608 <= _2597;
        else
            _2608 <= _2606;
    end
    assign _4848 = _2608 == _2605;
    assign _4849 = _4848 ? _4823 : _4847;
    assign _3355 = _4849;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3357 <= _3354;
        else
            _3357 <= _3355;
    end
    assign _5255 = _3357 & _3349;
    assign _5256 = _5255 ? _3385 : _3372;

    /* aliases */

    /* output assignments */
    assign next_pc = _5256;
    assign reg_op1 = _2664;
    assign reg_op2 = _2660;
    assign trap = _2656;
    assign mem_do_rinst = _2652;
    assign mem_do_wdata = _2648;
    assign mem_do_rdata = _2644;
    assign mem_wordsize = _2640;
    assign mem_do_prefetch = _2636;
    assign pcpi_valid = _2632;
    assign decoder_trigger = _2628;
    assign decoder_trigger_q = _2624;
    assign decoder_pseudo_trigger = _2620;
    assign eoi = _2616;
    assign ascii_state = ascii_state_0;

endmodule
