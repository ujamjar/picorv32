module opicorv32_rv32 (
    pcpi_rd,
    pcpi_wait,
    irq,
    pcpi_wr,
    pcpi_ready,
    mem_rdata,
    resetn,
    clk,
    mem_ready,
    trap,
    mem_valid,
    mem_instr,
    mem_addr,
    mem_wdata,
    mem_wstrb,
    mem_la_read,
    mem_la_write,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    pcpi_valid,
    pcpi_insn,
    pcpi_rs1,
    pcpi_rs2,
    eoi
);

    input [31:0] pcpi_rd;
    input pcpi_wait;
    input [31:0] irq;
    input pcpi_wr;
    input pcpi_ready;
    input [31:0] mem_rdata;
    input resetn;
    input clk;
    input mem_ready;
    output trap;
    output mem_valid;
    output mem_instr;
    output [31:0] mem_addr;
    output [31:0] mem_wdata;
    output [3:0] mem_wstrb;
    output mem_la_read;
    output mem_la_write;
    output [31:0] mem_la_addr;
    output [31:0] mem_la_wdata;
    output [3:0] mem_la_wstrb;
    output pcpi_valid;
    output [31:0] pcpi_insn;
    output [31:0] pcpi_rs1;
    output [31:0] pcpi_rs2;
    output [31:0] eoi;

    /* signal declarations */
    wire [31:0] _6750 = 32'b00000000000000000000000000000000;
    wire [31:0] _6748 = 32'b00000000000000000000000000000000;
    wire [31:0] _7799;
    wire [31:0] _7800;
    wire [31:0] _9325;
    wire [31:0] _9326;
    wire [31:0] _9327;
    wire [31:0] _9328;
    wire [31:0] _7878 = 32'b00000000000000000000000000000000;
    wire [31:0] _9329;
    wire [31:0] _9330;
    wire [31:0] _9331;
    wire [31:0] _9332;
    wire [31:0] _9333;
    wire [31:0] _9334;
    wire _9335;
    wire [31:0] _9336;
    wire _9337;
    wire [31:0] _9338;
    wire [31:0] _6749;
    reg [31:0] _6751;
    wire [31:0] _5661;
    wire [3:0] _5646;
    wire [31:0] _5647;
    wire [31:0] _5648;
    wire _6587;
    wire _6588;
    wire _5649;
    wire _6589;
    wire _6590;
    wire _6571;
    wire _6591;
    wire _6592;
    wire _5650;
    wire [3:0] _6687 = 4'b0000;
    wire [3:0] _6685 = 4'b0000;
    wire [3:0] _6693 = 4'b0000;
    wire [3:0] _6617 = 4'b1000;
    wire [3:0] _6616 = 4'b0100;
    wire [3:0] _6615 = 4'b0010;
    wire [3:0] _6614 = 4'b0001;
    wire [1:0] _6618;
    reg [3:0] _6619;
    wire [3:0] _6621 = 4'b1100;
    wire [3:0] _6620 = 4'b0011;
    wire _6622;
    wire [3:0] _6623;
    wire [3:0] _6624 = 4'b1111;
    reg [3:0] _6625;
    wire [3:0] _6701;
    wire _6702;
    wire [3:0] _6703;
    wire [3:0] _6686;
    reg [3:0] _6688;
    wire [3:0] _5654;
    wire [31:0] _6683 = 32'b00000000000000000000000000000000;
    wire [31:0] _6681 = 32'b00000000000000000000000000000000;
    wire [7:0] _6609;
    wire [15:0] _6610;
    wire [31:0] _6611;
    wire [15:0] _6606;
    wire [31:0] _6607;
    reg [31:0] _6613;
    wire _6704;
    wire [31:0] _6705;
    wire [31:0] _6682;
    reg [31:0] _6684;
    wire [31:0] _5655;
    wire [31:0] _6679 = 32'b00000000000000000000000000000000;
    wire [31:0] _6677 = 32'b00000000000000000000000000000000;
    wire _9390;
    wire [31:0] _9391;
    wire [31:0] _5674;
    wire [1:0] _6593 = 2'b00;
    wire [29:0] _6594;
    wire [31:0] _6595;
    wire _6596;
    wire [31:0] _6597;
    wire _6706;
    wire [31:0] _6707;
    wire [31:0] _6678;
    reg [31:0] _6680;
    wire [31:0] _5656;
    wire _6690 = 1'b0;
    wire _6694;
    wire _6697;
    wire _6698;
    wire _6699;
    wire _6700;
    wire _6689;
    reg _6691;
    wire _5657;
    wire _5658;
    wire _6790 = 1'b0;
    wire _6788 = 1'b0;
    wire _8267 = 1'b0;
    wire [2:0] _6742 = 3'b000;
    wire [2:0] _6732 = 3'b000;
    wire [2:0] _9339;
    wire [2:0] _9340;
    wire [2:0] _9341;
    wire [2:0] _9342;
    wire [2:0] _9343;
    wire [2:0] _9344;
    wire [2:0] _9345;
    wire [2:0] _9346;
    wire [2:0] _9347;
    wire [2:0] _9348;
    wire [2:0] _9349;
    wire [2:0] _9350;
    wire [2:0] _9351;
    wire [2:0] _9352;
    wire [2:0] _9353;
    wire [2:0] _9354;
    wire [2:0] _9355;
    wire [2:0] _9356;
    wire [2:0] _9357;
    wire [2:0] _9358;
    wire [2:0] _9359;
    wire [2:0] _9360;
    wire [2:0] _9361;
    wire [2:0] _9362;
    wire [2:0] _6739 = 3'b001;
    wire [2:0] _9363;
    wire [2:0] _9364;
    wire [2:0] _9365;
    wire [2:0] _9366;
    wire [2:0] _9367;
    wire [2:0] _9368;
    wire [2:0] _9369;
    wire [2:0] _9370;
    wire [2:0] _9371;
    wire [2:0] _9372;
    wire [2:0] _9373;
    wire [2:0] _9374;
    wire _6770 = 1'b0;
    wire _6768 = 1'b0;
    wire _8080 = 1'b0;
    wire _7674;
    wire _7675;
    wire _7676;
    wire _7677;
    wire _7678;
    wire _9288;
    wire _9289;
    wire _9290;
    wire _9291;
    wire _9292;
    wire _9293;
    wire _6572;
    wire _6581;
    wire _6582;
    wire _6583;
    wire [1:0] _6569 = 2'b00;
    wire [1:0] _6563 = 2'b00;
    wire [1:0] _6718;
    wire [1:0] _6719;
    wire _6692;
    wire [1:0] _6720;
    wire [1:0] _6721;
    wire [1:0] _6722;
    wire _6786 = 1'b0;
    wire _6784 = 1'b0;
    wire _8076 = 1'b1;
    wire _8079 = 1'b0;
    wire _7689 = 1'b1;
    wire _9174;
    wire _9175;
    wire _9176;
    wire _9177;
    wire _9178;
    wire _9179;
    wire _9180;
    wire _9181;
    wire _9182;
    wire _9183;
    wire _9184;
    wire _9185;
    wire _9186;
    wire _9187;
    wire _9188;
    wire _9189;
    wire _9190;
    wire _9191;
    wire _9192;
    wire _9193;
    wire _9194;
    wire _9195;
    wire _9196;
    wire _9197;
    wire _9198;
    wire _9199;
    wire _9200;
    wire _9201;
    wire _9202;
    wire _9203;
    wire _9204;
    wire _9205;
    wire _9206;
    wire _9207;
    wire _9208;
    wire _9209;
    wire _9210;
    wire _9211;
    wire _9212;
    wire _9213;
    wire _9214;
    wire _9215;
    wire _9216;
    wire _9217;
    wire _9218;
    wire _9219;
    wire _9220;
    wire _9221;
    wire _9222;
    wire _9223;
    wire _9224;
    wire _9225;
    wire _9226;
    wire _9227;
    wire _9228;
    wire _9229;
    wire _9230;
    wire _9231;
    wire _9232;
    wire _9233;
    wire _9234;
    wire _9235;
    wire _9236;
    wire _9237;
    wire _7682 = 1'b1;
    wire _7679 = 1'b0;
    wire _9238;
    wire _7803 = 1'b1;
    wire _7813;
    wire _7814;
    wire _7815;
    wire _9171;
    wire _9172;
    wire _9173;
    wire _9239;
    wire _9240;
    wire _9241;
    wire _7922 = 1'b1;
    wire _9242;
    wire _9243;
    wire _9244;
    wire _7833 = 1'b1;
    wire _7827 = 1'b1;
    wire _7826;
    wire _9245;
    wire _7828;
    wire _9246;
    wire _9247;
    wire _9248;
    wire _9249;
    wire _9250;
    wire _9251;
    wire _9252;
    wire _9253;
    wire _9254;
    wire _9255;
    wire _9256;
    wire _9257;
    wire _9258;
    wire _7937 = 1'b1;
    wire _9259;
    wire _7929 = 1'b1;
    wire _7928;
    wire _9260;
    wire _7930;
    wire _9261;
    wire _9262;
    wire _9263;
    wire _9264;
    wire _9265;
    wire _9266;
    wire _9267;
    wire _9268;
    wire _9269;
    wire _9270;
    wire _9271;
    wire _9272;
    wire _7945 = 1'b1;
    wire _8279;
    wire _6444 = 1'b0;
    wire _6441;
    wire _6440;
    wire _6439;
    wire _6442;
    wire _6443;
    reg is_lui_auipc_jal;
    wire _6393 = 1'b0;
    wire [6:0] _6370 = 7'b0100000;
    wire [6:0] _6369;
    wire _6371;
    wire [2:0] _6373 = 3'b101;
    wire [2:0] _6372;
    wire _6374;
    wire _6375;
    wire [6:0] _6377 = 7'b0000000;
    wire [6:0] _6376;
    wire _6378;
    wire [2:0] _6380 = 3'b101;
    wire [2:0] _6379;
    wire _6381;
    wire _6382;
    wire [6:0] _6384 = 7'b0000000;
    wire [6:0] _6383;
    wire _6385;
    wire [2:0] _6387 = 3'b001;
    wire [2:0] _6386;
    wire _6388;
    wire _6389;
    wire _6390;
    wire _6391;
    wire _6392;
    reg is_slli_srli_srai;
    wire _6367 = 1'b0;
    wire [2:0] _6343 = 3'b111;
    wire [2:0] _6342;
    wire _6344;
    wire [2:0] _6346 = 3'b110;
    wire [2:0] _6345;
    wire _6347;
    wire [2:0] _6349 = 3'b100;
    wire [2:0] _6348;
    wire _6350;
    wire [2:0] _6352 = 3'b011;
    wire [2:0] _6351;
    wire _6353;
    wire [2:0] _6355 = 3'b010;
    wire [2:0] _6354;
    wire _6356;
    wire [2:0] _6358 = 3'b000;
    wire [2:0] _6357;
    wire _6359;
    wire _6360;
    wire _6361;
    wire _6362;
    wire _6363;
    wire _6364;
    wire _6365;
    wire _6366;
    reg is_jalr_addi_slti_sltiu_xori_ori_andi;
    wire _6340 = 1'b0;
    wire [6:0] _6317 = 7'b0100000;
    wire [6:0] _6316;
    wire _6318;
    wire [2:0] _6320 = 3'b101;
    wire [2:0] _6319;
    wire _6321;
    wire _6322;
    wire [6:0] _6324 = 7'b0000000;
    wire [6:0] _6323;
    wire _6325;
    wire [2:0] _6327 = 3'b101;
    wire [2:0] _6326;
    wire _6328;
    wire _6329;
    wire [6:0] _6331 = 7'b0000000;
    wire [6:0] _6330;
    wire _6332;
    wire [2:0] _6334 = 3'b001;
    wire [2:0] _6333;
    wire _6335;
    wire _6336;
    wire _6337;
    wire _6338;
    wire _6339;
    reg is_sll_srl_sra;
    wire _6437 = 1'b0;
    wire _6431;
    wire _6430;
    wire _6429;
    wire _6428;
    wire _6427;
    wire _6426;
    wire _6432;
    wire _6433;
    wire _6434;
    wire _6435;
    wire _6436;
    reg is_lui_auipc_jal_jalr_addi_add;
    wire _6424 = 1'b0;
    wire _6421;
    wire _6420;
    wire _6419;
    wire _6422;
    wire _6423;
    reg is_slti_blt_slt;
    wire _6417 = 1'b0;
    wire _6414;
    wire _6413;
    wire _6412;
    wire _6415;
    wire _6416;
    reg is_sltiu_bltu_sltu;
    wire _6410 = 1'b0;
    wire _6407;
    wire _6406;
    wire _6405;
    wire _6408;
    wire _6409;
    reg is_lbu_lhu_lw;
    wire _6403 = 1'b0;
    wire _6398;
    wire _6397;
    wire _6396;
    wire _6395;
    wire _6399;
    wire _6400;
    wire _6401;
    wire _6402;
    reg is_compare;
    wire _6312;
    wire _6311;
    wire _6310;
    wire _5901 = 1'b0;
    wire [6:0] _5893 = 7'b0000101;
    wire [6:0] _5892;
    wire _5894;
    wire [6:0] _5896 = 7'b0001011;
    wire [6:0] _5895;
    wire _5897;
    wire _5898;
    wire _5899;
    wire _5900;
    reg instr_timer;
    wire _5911 = 1'b0;
    wire [6:0] _5904 = 7'b0000011;
    wire [6:0] _5903;
    wire _5905;
    wire [6:0] _5907 = 7'b0001011;
    wire [6:0] _5906;
    wire _5908;
    wire _5909;
    wire _5910;
    reg instr_maskirq;
    wire _5922 = 1'b0;
    wire [6:0] _5914 = 7'b0000001;
    wire [6:0] _5913;
    wire _5915;
    wire [6:0] _5917 = 7'b0001011;
    wire [6:0] _5916;
    wire _5918;
    wire _5919;
    wire _5920;
    wire _5921;
    reg instr_setq;
    wire _5933 = 1'b0;
    wire [6:0] _5925 = 7'b0000000;
    wire [6:0] _5924;
    wire _5926;
    wire [6:0] _5928 = 7'b0001011;
    wire [6:0] _5927;
    wire _5929;
    wire _5930;
    wire _5931;
    wire _5932;
    reg instr_getq;
    wire _5943 = 1'b0;
    wire [19:0] _5936 = 20'b11001000001000000010;
    wire [19:0] _5935;
    wire _5937;
    wire [6:0] _5939 = 7'b1110011;
    wire [6:0] _5938;
    wire _5940;
    wire _5941;
    wire _5942;
    reg instr_rdinstrh;
    wire _5953 = 1'b0;
    wire [19:0] _5946 = 20'b11000000001000000010;
    wire [19:0] _5945;
    wire _5947;
    wire [6:0] _5949 = 7'b1110011;
    wire [6:0] _5948;
    wire _5950;
    wire _5951;
    wire _5952;
    reg instr_rdinstr;
    wire _5971 = 1'b0;
    wire [19:0] _5956 = 20'b11001000000100000010;
    wire [19:0] _5955;
    wire _5957;
    wire [6:0] _5959 = 7'b1110011;
    wire [6:0] _5958;
    wire _5960;
    wire _5961;
    wire [19:0] _5963 = 20'b11001000000000000010;
    wire [19:0] _5962;
    wire _5964;
    wire [6:0] _5966 = 7'b1110011;
    wire [6:0] _5965;
    wire _5967;
    wire _5968;
    wire _5969;
    wire _5970;
    reg instr_rdcycleh;
    wire _5989 = 1'b0;
    wire [19:0] _5974 = 20'b11000000000100000010;
    wire [19:0] _5973;
    wire _5975;
    wire [6:0] _5977 = 7'b1110011;
    wire [6:0] _5976;
    wire _5978;
    wire _5979;
    wire [19:0] _5981 = 20'b11000000000000000010;
    wire [19:0] _5980;
    wire _5982;
    wire [6:0] _5984 = 7'b1110011;
    wire [6:0] _5983;
    wire _5985;
    wire _5986;
    wire _5987;
    wire _5988;
    reg instr_rdcycle;
    wire _5999 = 1'b0;
    wire [6:0] _5992 = 7'b0000000;
    wire [6:0] _5991;
    wire _5993;
    wire [2:0] _5995 = 3'b111;
    wire [2:0] _5994;
    wire _5996;
    wire _5997;
    wire _5998;
    reg instr_and;
    wire _6009 = 1'b0;
    wire [6:0] _6002 = 7'b0000000;
    wire [6:0] _6001;
    wire _6003;
    wire [2:0] _6005 = 3'b110;
    wire [2:0] _6004;
    wire _6006;
    wire _6007;
    wire _6008;
    reg instr_or;
    wire _6019 = 1'b0;
    wire [6:0] _6012 = 7'b0100000;
    wire [6:0] _6011;
    wire _6013;
    wire [2:0] _6015 = 3'b101;
    wire [2:0] _6014;
    wire _6016;
    wire _6017;
    wire _6018;
    reg instr_sra;
    wire _6029 = 1'b0;
    wire [6:0] _6022 = 7'b0000000;
    wire [6:0] _6021;
    wire _6023;
    wire [2:0] _6025 = 3'b101;
    wire [2:0] _6024;
    wire _6026;
    wire _6027;
    wire _6028;
    reg instr_srl;
    wire _6039 = 1'b0;
    wire [6:0] _6032 = 7'b0000000;
    wire [6:0] _6031;
    wire _6033;
    wire [2:0] _6035 = 3'b100;
    wire [2:0] _6034;
    wire _6036;
    wire _6037;
    wire _6038;
    reg instr_xor;
    wire _6049 = 1'b0;
    wire [6:0] _6042 = 7'b0000000;
    wire [6:0] _6041;
    wire _6043;
    wire [2:0] _6045 = 3'b011;
    wire [2:0] _6044;
    wire _6046;
    wire _6047;
    wire _6048;
    reg instr_sltu;
    wire _6059 = 1'b0;
    wire [6:0] _6052 = 7'b0000000;
    wire [6:0] _6051;
    wire _6053;
    wire [2:0] _6055 = 3'b010;
    wire [2:0] _6054;
    wire _6056;
    wire _6057;
    wire _6058;
    reg instr_slt;
    wire _6069 = 1'b0;
    wire [6:0] _6062 = 7'b0000000;
    wire [6:0] _6061;
    wire _6063;
    wire [2:0] _6065 = 3'b001;
    wire [2:0] _6064;
    wire _6066;
    wire _6067;
    wire _6068;
    reg instr_sll;
    wire _6079 = 1'b0;
    wire [6:0] _6072 = 7'b0100000;
    wire [6:0] _6071;
    wire _6073;
    wire [2:0] _6075 = 3'b000;
    wire [2:0] _6074;
    wire _6076;
    wire _6077;
    wire _6078;
    reg instr_sub;
    wire _6089 = 1'b0;
    wire [6:0] _6082 = 7'b0000000;
    wire [6:0] _6081;
    wire _6083;
    wire [2:0] _6085 = 3'b000;
    wire [2:0] _6084;
    wire _6086;
    wire _5890 = 1'b0;
    wire [6:0] _5888 = 7'b0110011;
    wire [6:0] _5887;
    wire _5889;
    reg is_alu_reg_reg;
    wire _6087;
    wire _6088;
    reg instr_add;
    wire _6099 = 1'b0;
    wire [6:0] _6092 = 7'b0100000;
    wire [6:0] _6091;
    wire _6093;
    wire [2:0] _6095 = 3'b101;
    wire [2:0] _6094;
    wire _6096;
    wire _6097;
    wire _6098;
    reg instr_srai;
    wire _6109 = 1'b0;
    wire [6:0] _6102 = 7'b0000000;
    wire [6:0] _6101;
    wire _6103;
    wire [2:0] _6105 = 3'b101;
    wire [2:0] _6104;
    wire _6106;
    wire _6107;
    wire _6108;
    reg instr_srli;
    wire _6119 = 1'b0;
    wire [6:0] _6112 = 7'b0000000;
    wire [6:0] _6111;
    wire _6113;
    wire [2:0] _6115 = 3'b001;
    wire [2:0] _6114;
    wire _6116;
    wire _6117;
    wire _6118;
    reg instr_slli;
    wire _6125 = 1'b0;
    wire [2:0] _6122 = 3'b111;
    wire [2:0] _6121;
    wire _6123;
    wire _6124;
    reg instr_andi;
    wire _6131 = 1'b0;
    wire [2:0] _6128 = 3'b110;
    wire [2:0] _6127;
    wire _6129;
    wire _6130;
    reg instr_ori;
    wire _6137 = 1'b0;
    wire [2:0] _6134 = 3'b100;
    wire [2:0] _6133;
    wire _6135;
    wire _6136;
    reg instr_xori;
    wire _6143 = 1'b0;
    wire [2:0] _6140 = 3'b011;
    wire [2:0] _6139;
    wire _6141;
    wire _6142;
    reg instr_sltiu;
    wire _6149 = 1'b0;
    wire [2:0] _6146 = 3'b010;
    wire [2:0] _6145;
    wire _6147;
    wire _6148;
    reg instr_slti;
    wire _6155 = 1'b0;
    wire [2:0] _6152 = 3'b000;
    wire [2:0] _6151;
    wire _6153;
    wire _5885 = 1'b0;
    wire [6:0] _5883 = 7'b0010011;
    wire [6:0] _5882;
    wire _5884;
    reg is_alu_reg_imm;
    wire _6154;
    reg instr_addi;
    wire _6161 = 1'b0;
    wire [2:0] _6158 = 3'b010;
    wire [2:0] _6157;
    wire _6159;
    wire _6160;
    reg instr_sw;
    wire _6167 = 1'b0;
    wire [2:0] _6164 = 3'b001;
    wire [2:0] _6163;
    wire _6165;
    wire _6166;
    reg instr_sh;
    wire _6173 = 1'b0;
    wire [2:0] _6170 = 3'b000;
    wire [2:0] _6169;
    wire _6171;
    wire _5880 = 1'b0;
    wire [6:0] _5878 = 7'b0100011;
    wire [6:0] _5877;
    wire _5879;
    reg is_sb_sh_sw;
    wire _6172;
    reg instr_sb;
    wire _6179 = 1'b0;
    wire [2:0] _6176 = 3'b101;
    wire [2:0] _6175;
    wire _6177;
    wire _6178;
    reg instr_lhu;
    wire _6185 = 1'b0;
    wire [2:0] _6182 = 3'b100;
    wire [2:0] _6181;
    wire _6183;
    wire _6184;
    reg instr_lbu;
    wire _6191 = 1'b0;
    wire [2:0] _6188 = 3'b010;
    wire [2:0] _6187;
    wire _6189;
    wire _6190;
    reg instr_lw;
    wire _6197 = 1'b0;
    wire [2:0] _6194 = 3'b001;
    wire [2:0] _6193;
    wire _6195;
    wire _6196;
    reg instr_lh;
    wire _6203 = 1'b0;
    wire [2:0] _6200 = 3'b000;
    wire [2:0] _6199;
    wire _6201;
    wire _5875 = 1'b0;
    wire [6:0] _5873 = 7'b0000011;
    wire [6:0] _5872;
    wire _5874;
    reg is_lb_lh_lw_lbu_lhu;
    wire _6202;
    reg instr_lb;
    wire _6209 = 1'b0;
    wire [2:0] _6206 = 3'b111;
    wire [2:0] _6205;
    wire _6207;
    wire _6208;
    reg instr_bgeu;
    wire _6215 = 1'b0;
    wire [2:0] _6212 = 3'b110;
    wire [2:0] _6211;
    wire _6213;
    wire _6214;
    reg instr_bltu;
    wire _6221 = 1'b0;
    wire [2:0] _6218 = 3'b101;
    wire [2:0] _6217;
    wire _6219;
    wire _6220;
    reg instr_bge;
    wire _6227 = 1'b0;
    wire [2:0] _6224 = 3'b100;
    wire [2:0] _6223;
    wire _6225;
    wire _6226;
    reg instr_blt;
    wire _6233 = 1'b0;
    wire [2:0] _6230 = 3'b001;
    wire [2:0] _6229;
    wire _6231;
    wire _6232;
    reg instr_bne;
    wire _5845;
    wire _6762 = 1'b0;
    wire _6760 = 1'b0;
    wire _7946 = 1'b0;
    wire _7412;
    wire _7409;
    wire _7410;
    wire _7418;
    wire [30:0] _7398;
    wire _7399;
    wire _7400;
    wire [31:0] _7401;
    wire [30:0] _7402;
    wire _7403;
    wire _7404;
    wire [31:0] _7405;
    wire _7406;
    wire _7407;
    wire _7395;
    wire _7396;
    wire _7416;
    wire _7420;
    wire [30:0] _7385;
    wire _7386;
    wire _7387;
    wire [31:0] _7388;
    wire [30:0] _7389;
    wire _7390;
    wire _7391;
    wire [31:0] _7392;
    wire _7393;
    wire [31:0] _6798 = 32'b00000000000000000000000000000000;
    wire [31:0] _6796 = 32'b00000000000000000000000000000000;
    wire [31:0] _9128;
    wire [31:0] _7891 = 32'b00000000000000000000000000000000;
    wire _7892;
    wire [31:0] _7893;
    wire [31:0] _7927 = 32'b00000000000000000000000000000000;
    wire [31:0] _9129;
    wire [31:0] _9130;
    wire [31:0] _9131;
    wire [31:0] _9132;
    wire [31:0] _9133;
    wire [31:0] _9134;
    wire [31:0] _9135;
    wire [31:0] _9136;
    wire [3:0] _7991 = 4'b0000;
    wire [27:0] _7992;
    wire [31:0] _7993;
    wire [27:0] _7985;
    wire [3:0] _7986 = 4'b0000;
    wire [31:0] _7987;
    wire [31:0] _7997;
    wire [27:0] _7976;
    wire _7977;
    wire [1:0] _7978;
    wire [3:0] _7979;
    wire [31:0] _7981;
    wire _7988;
    wire _7989;
    wire _7990;
    wire _7994;
    wire _7995;
    wire _7996;
    wire _7998;
    wire [31:0] _7999;
    wire _7964 = 1'b0;
    wire [30:0] _7965;
    wire [31:0] _7966;
    wire [30:0] _7958;
    wire _7959 = 1'b0;
    wire [31:0] _7960;
    wire [31:0] _7970;
    wire [30:0] _7952;
    wire _7953;
    wire [31:0] _7954;
    wire _7961;
    wire _7962;
    wire _7963;
    wire _7967;
    wire _7968;
    wire _7969;
    wire _7971;
    wire [31:0] _7972;
    wire [31:0] _9137;
    wire [4:0] _8004 = 5'b00000;
    wire [4:0] _7523 = 5'b00000;
    wire [4:0] _7521 = 5'b00000;
    wire [4:0] _7923;
    wire [4:0] _8682;
    wire [4:0] _8683;
    wire [4:0] _7831;
    wire [4:0] _7829;
    wire [4:0] _8684;
    wire [4:0] _8685;
    wire [4:0] _8686;
    wire [4:0] _8687;
    wire [4:0] _8688;
    wire [4:0] _8689;
    wire [4:0] _8690;
    wire [4:0] _8691;
    wire [4:0] _8692;
    wire [4:0] _8693;
    wire [4:0] _8694;
    wire [4:0] _8695;
    wire _7201;
    wire _7202;
    wire [31:0] _7204 = 32'b00000000000000000000000000000000;
    wire [31:0] _7203 = 32'b00000000000000000000000000000000;
    wire [31:0] _7808 = 32'b00000000000000000000000000000100;
    wire [31:0] _7809;
    wire [31:0] _9103;
    wire [31:0] _7807;
    wire [31:0] _9104;
    wire [31:0] _7506 = 32'b00000000000000000000000000000000;
    wire [31:0] _7690 = 32'b00000000000000000000000000000100;
    wire [31:0] _7691;
    wire _8805;
    wire _8806;
    wire _8807;
    wire _8808;
    wire _8809;
    wire _8810;
    wire _8811;
    wire _8812;
    wire _8813;
    wire _8814;
    wire _8815;
    wire _8816;
    wire _8817;
    wire _8818;
    wire _8819;
    wire _8820;
    wire _8821;
    wire _8822;
    wire _8823;
    wire _8824;
    wire _8825;
    wire _8826;
    wire _8827;
    wire _8828;
    wire _8829;
    wire _8830;
    wire _8831;
    wire _8832;
    wire _8833;
    wire _8834;
    wire _8835;
    wire _8836;
    wire _8837;
    wire _8838;
    wire _8839;
    wire _8840;
    wire _8841;
    wire _8842;
    wire _8843;
    wire _8844;
    wire _8845;
    wire _8846;
    wire _8847;
    wire _8848;
    wire _8849;
    wire _8850;
    wire _8851;
    wire _8852;
    wire _8853;
    wire _8854;
    wire _8855;
    wire _8856;
    wire _8857;
    wire _8858;
    wire _8859;
    wire _8860;
    wire _8861;
    wire _8862;
    wire _8863;
    wire _8864;
    wire _8865;
    wire _8866;
    wire _8867;
    wire [31:0] _8868;
    wire [31:0] _5638;
    wire [31:0] _7681;
    wire [31:0] _7686 = 32'b00000000000000000000000000000100;
    wire [31:0] _7687;
    wire [31:0] _8869;
    wire [31:0] _7515 = 32'b00000000000000000000000000000000;
    wire [31:0] _7513 = 32'b00000000000000000000000000000000;
    wire [31:0] _7449;
    wire [31:0] _7447;
    wire [31:0] _7455;
    wire [30:0] _7443 = 31'b0000000000000000000000000000000;
    wire [31:0] _7445;
    wire [31:0] _7432;
    wire [31:0] _7453;
    wire [31:0] _7457;
    wire [31:0] _7428;
    wire [31:0] _7424;
    wire _7429;
    wire _7430;
    wire _7431;
    wire [31:0] _7451;
    wire _7433;
    wire _7434;
    wire _7435;
    wire _7446;
    wire _7454;
    wire _7448;
    wire _7450;
    wire _7456;
    wire _7458;
    wire [31:0] _7459;
    wire [31:0] _7514;
    reg [31:0] _7516;
    wire [31:0] _7519 = 32'b00000000000000000000000000000000;
    wire [31:0] _7517 = 32'b00000000000000000000000000000000;
    wire _8704;
    wire _8705;
    wire _8706;
    wire _8707;
    wire _8708;
    wire _8709;
    wire _8710;
    wire _8711;
    wire _8712;
    wire _8713;
    wire _8714;
    wire _8715;
    wire _8716;
    wire _8717;
    wire _8718;
    wire _8719;
    wire _8720;
    wire _8721;
    wire _8722;
    wire _8723;
    wire _8724;
    wire _8725;
    wire _8726;
    wire _8727;
    wire _8728;
    wire _8729;
    wire _8730;
    wire _8731;
    wire _8732;
    wire _8733;
    wire _8734;
    wire _8735;
    wire _8736;
    wire _8737;
    wire _8738;
    wire _8739;
    wire _8740;
    wire _8741;
    wire _8742;
    wire _8743;
    wire _8744;
    wire _8745;
    wire _8746;
    wire _8747;
    wire _8748;
    wire _8749;
    wire _8750;
    wire _8751;
    wire _8752;
    wire _8753;
    wire _8754;
    wire _8755;
    wire _8756;
    wire _8757;
    wire _8758;
    wire _8759;
    wire _8760;
    wire _8761;
    wire _8762;
    wire _8763;
    wire _8764;
    wire _8765;
    wire _8766;
    wire [31:0] _8767;
    wire [31:0] _8768;
    wire [31:0] _8769;
    wire [31:0] _8770;
    wire [31:0] _8771;
    wire [31:0] _8772;
    wire [31:0] _7902;
    wire [63:0] _7479 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7477 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _8096 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _8097;
    wire [63:0] _9007;
    wire [63:0] _7478;
    reg [63:0] count_cycle;
    wire [31:0] _7900;
    wire [31:0] _7906;
    wire [31:0] _7898;
    wire [63:0] _7475 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7473 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7684 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _7685;
    wire [63:0] _9008;
    wire [63:0] _9009;
    wire [63:0] _9010;
    wire [63:0] _9011;
    wire _9012;
    wire [63:0] _9013;
    wire [63:0] _7474;
    reg [63:0] _7476;
    wire [31:0] _7896;
    wire _7899;
    wire [31:0] _7904;
    wire _7901;
    wire _7903;
    wire _7907;
    wire [31:0] _7908;
    wire [31:0] _8773;
    wire [31:0] _8774;
    wire [31:0] _8775;
    wire [31:0] _8776;
    wire [31:0] _8777;
    wire [31:0] _8778;
    wire [31:0] _8779;
    wire [31:0] _8780;
    wire [31:0] _5828 = 32'b00000000000000000000000000000000;
    wire [31:0] _5827 = 32'b00000000000000000000000000000000;
    wire [31:0] _5825;
    wire [63:0] _5738 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5736 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5778 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5741;
    wire [63:0] _5734 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5732 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5777 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5751 = 1'b0;
    wire [63:0] _5745;
    wire [63:0] _5726 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5724 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5786;
    wire [1:0] _5787;
    wire [3:0] _5788;
    wire [7:0] _5789;
    wire [15:0] _5790;
    wire [31:0] _5791;
    wire [63:0] _5793;
    wire [31:0] _6794 = 32'b00000000000000000000000000000000;
    wire [31:0] _6792 = 32'b00000000000000000000000000000000;
    wire [31:0] _9151;
    wire [31:0] _9152;
    wire [31:0] _7926 = 32'b00000000000000000000000000000000;
    wire [31:0] _9153;
    wire _7830;
    wire [31:0] _9154;
    wire _7832;
    wire [31:0] _9155;
    wire _7834;
    wire [31:0] _9156;
    wire [31:0] _9157;
    wire [31:0] _9158;
    wire [31:0] _9159;
    wire [31:0] _9160;
    wire [31:0] _9161;
    wire [31:0] _9162;
    wire [31:0] _9163;
    wire [31:0] _9164;
    wire _9165;
    wire [31:0] _9166;
    wire _9167;
    wire [31:0] _9168;
    wire [31:0] _6793;
    reg [31:0] _6795;
    wire [31:0] _5672;
    wire [31:0] _5783 = 32'b00000000000000000000000000000000;
    wire [63:0] _5785;
    wire [63:0] _5794;
    wire _5757 = 1'b0;
    wire [62:0] _5758;
    wire [63:0] _5759;
    wire [63:0] _5819;
    wire [63:0] _5725;
    reg [63:0] _5727;
    wire [63:0] _5746;
    wire [63:0] _5747;
    wire [63:0] _5748;
    wire [63:0] _5744;
    wire _5749;
    wire [63:0] _5750;
    wire [62:0] _5752;
    wire [63:0] _5753;
    wire [63:0] _5817;
    wire [63:0] _5733;
    reg [63:0] _5735;
    wire [63:0] _5740;
    wire [63:0] _5730 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5728 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5802;
    wire [1:0] _5803;
    wire [3:0] _5804;
    wire [7:0] _5805;
    wire [15:0] _5806;
    wire [31:0] _5807;
    wire [63:0] _5809;
    wire [31:0] _5799 = 32'b00000000000000000000000000000000;
    wire [63:0] _5801;
    wire _5717;
    wire [63:0] _5810;
    wire [62:0] _5754;
    wire _5755 = 1'b0;
    wire [63:0] _5756;
    wire [63:0] _5818;
    wire [63:0] _5729;
    reg [63:0] _5731;
    wire _5742;
    wire [63:0] _5743;
    wire [63:0] _5816;
    wire [63:0] _5737;
    reg [63:0] _5739;
    wire [31:0] _5824;
    wire [31:0] _5826;
    reg [31:0] _5829;
    wire [31:0] _5838 = 32'b00000000000000000000000000000000;
    wire [31:0] _5839;
    wire [31:0] _5840;
    wire [31:0] _5636;
    wire [31:0] _8781;
    wire [31:0] _8782;
    wire [31:0] _7509 = 32'b00000000000000000000000000000000;
    wire [31:0] _39 = 32'b00000000000000000000000000000000;
    wire _8803;
    wire [31:0] _8804;
    wire [31:0] _7508;
    reg [31:0] _7510;
    wire [31:0] _7949;
    wire [31:0] _8783;
    wire [15:0] _8037;
    wire _8038;
    wire [1:0] _8039;
    wire [3:0] _8040;
    wire [7:0] _8041;
    wire [15:0] _8042;
    wire [31:0] _8044;
    wire [31:0] _8045;
    wire [7:0] _6650;
    wire [23:0] _6655 = 24'b000000000000000000000000;
    wire [31:0] _6657;
    wire [7:0] _6642;
    wire [23:0] _6647 = 24'b000000000000000000000000;
    wire [31:0] _6649;
    wire [7:0] _6634;
    wire [23:0] _6639 = 24'b000000000000000000000000;
    wire [31:0] _6641;
    wire [7:0] _6626;
    wire [23:0] _6631 = 24'b000000000000000000000000;
    wire [31:0] _6633;
    wire [1:0] _6658;
    reg [31:0] _6659;
    wire [15:0] _6660;
    wire [15:0] _6664 = 16'b0000000000000000;
    wire [31:0] _6666;
    wire [15:0] _6667;
    wire [15:0] _6671 = 16'b0000000000000000;
    wire [31:0] _6673;
    wire [31:0] _5673;
    wire _6674;
    wire [31:0] _6675;
    wire [1:0] _6774 = 2'b00;
    wire [1:0] _6772 = 2'b00;
    wire [1:0] _7812 = 2'b00;
    wire [1:0] _8017 = 2'b10;
    wire [1:0] _8015 = 2'b01;
    wire [1:0] _8019;
    wire [1:0] _8013 = 2'b00;
    wire _8016;
    wire _8018;
    wire _8020;
    wire [1:0] _8021;
    wire [1:0] _9278;
    wire [1:0] _9279;
    wire [1:0] _8062 = 2'b10;
    wire [1:0] _8058 = 2'b01;
    wire [1:0] _8066;
    wire [1:0] _8056 = 2'b00;
    wire _8059;
    wire _8060;
    wire _8061;
    wire _8063;
    wire _8064;
    wire _8065;
    wire _8067;
    wire [1:0] _8068;
    wire [1:0] _9280;
    wire [1:0] _9281;
    wire _9282;
    wire [1:0] _9283;
    wire _9284;
    wire [1:0] _9285;
    wire _9286;
    wire [1:0] _9287;
    wire [1:0] _6773;
    reg [1:0] _6775;
    wire [1:0] _5667;
    reg [31:0] _6676;
    wire [31:0] _5651;
    wire [7:0] _8028;
    wire _8029;
    wire [1:0] _8030;
    wire [3:0] _8031;
    wire [7:0] _8032;
    wire [15:0] _8033;
    wire [23:0] _8034;
    wire [31:0] _8036;
    wire _7499 = 1'b0;
    wire _7497 = 1'b0;
    wire _7791 = 1'b0;
    wire _8054;
    wire _8881;
    wire _8882;
    wire _8883;
    wire _8884;
    wire _8885;
    wire _8886;
    wire _7498;
    reg _7500;
    wire _7503 = 1'b0;
    wire _7501 = 1'b0;
    wire _7792 = 1'b0;
    wire _8055;
    wire _8875;
    wire _8876;
    wire _8877;
    wire _8878;
    wire _8879;
    wire _8880;
    wire _7502;
    reg _7504;
    wire _8046;
    wire [31:0] _8047;
    wire [31:0] _8784;
    wire [31:0] _8785;
    wire [31:0] _8265 = 32'b00000000000000000000000000000000;
    wire _8786;
    wire [31:0] _8787;
    wire _8788;
    wire [31:0] _8789;
    wire _8790;
    wire [31:0] _8791;
    wire _8792;
    wire [31:0] _8793;
    wire _8794;
    wire [31:0] _8795;
    wire _8796;
    wire [31:0] _8797;
    wire [31:0] _7518;
    reg [31:0] _7520;
    wire _7487 = 1'b0;
    wire _7485 = 1'b0;
    wire _7794 = 1'b0;
    wire _7942 = 1'b1;
    wire _8985;
    wire _8986;
    wire _8987;
    wire _8988;
    wire _8989;
    wire _7486;
    reg _7488;
    wire [31:0] _7810;
    wire [31:0] _7811;
    wire [31:0] _40 = 32'b00000000000000000000000000010000;
    wire [31:0] _8798;
    wire [31:0] _8799;
    wire [31:0] _8800;
    wire [31:0] _7511 = 32'b00000000000000000000000000000000;
    wire _8801;
    wire [31:0] _8802;
    wire [31:0] _7512;
    wire [31:0] _8870;
    wire [31:0] _8871;
    wire [31:0] _8872;
    wire _8873;
    wire [31:0] _8874;
    wire [31:0] _7505;
    reg [31:0] _7507;
    wire [31:0] _9105;
    wire [31:0] _7797;
    wire [31:0] _7798;
    wire [31:0] _9106;
    wire [31:0] _9107;
    wire [31:0] _9108;
    wire [31:0] _9109;
    wire _7483 = 1'b0;
    wire _7481 = 1'b0;
    wire _7680 = 1'b1;
    wire _7683;
    wire _8990;
    wire _7793 = 1'b0;
    wire _8991;
    wire _8992;
    wire _7717;
    wire _7718;
    wire _7719;
    wire _7722;
    wire _7723;
    wire _7724;
    wire _7725;
    wire _7726;
    wire _7727;
    wire _7728;
    wire _7729;
    wire _7730;
    wire _7731;
    wire _7732;
    wire _7733;
    wire _7734;
    wire _7735;
    wire _7736;
    wire _7737;
    wire _7738;
    wire _7739;
    wire _7740;
    wire _7741;
    wire _7742;
    wire _7743;
    wire _7744;
    wire _7745;
    wire _7746;
    wire _7747;
    wire _7748;
    wire _7749;
    wire _7750;
    wire _7751;
    wire _7752;
    wire [31:0] _7720;
    wire [31:0] _7721;
    wire _7753;
    wire _7754;
    wire _7755;
    wire _7756;
    wire _7757;
    wire _7758;
    wire _7759;
    wire _7760;
    wire _7761;
    wire _7762;
    wire _7763;
    wire _7764;
    wire _7765;
    wire _7766;
    wire _7767;
    wire _7768;
    wire _7769;
    wire _7770;
    wire _7771;
    wire _7772;
    wire _7773;
    wire _7774;
    wire _7775;
    wire _7776;
    wire _7777;
    wire _7778;
    wire _7779;
    wire _7780;
    wire _7781;
    wire _7782;
    wire _7783;
    wire _7784;
    wire _7531 = 1'b0;
    wire _7529 = 1'b0;
    wire _7804 = 1'b1;
    wire _8666;
    wire _7491 = 1'b0;
    wire _7489 = 1'b0;
    wire _7692 = 1'b1;
    wire _8893;
    wire _8894;
    wire _8895;
    wire _8896;
    wire _8897;
    wire _8898;
    wire _8899;
    wire _8900;
    wire _8901;
    wire _8902;
    wire _8903;
    wire _8904;
    wire _8905;
    wire _8906;
    wire _8907;
    wire _8908;
    wire _8909;
    wire _8910;
    wire _8911;
    wire _8912;
    wire _8913;
    wire _8914;
    wire _8915;
    wire _8916;
    wire _8917;
    wire _8918;
    wire _8919;
    wire _8920;
    wire _8921;
    wire _8922;
    wire _8923;
    wire _8924;
    wire _8925;
    wire _8926;
    wire _8927;
    wire _8928;
    wire _8929;
    wire _8930;
    wire _8931;
    wire _8932;
    wire _8933;
    wire _8934;
    wire _8935;
    wire _8936;
    wire _8937;
    wire _8938;
    wire _8939;
    wire _8940;
    wire _8941;
    wire _8942;
    wire _8943;
    wire _8944;
    wire _8945;
    wire _8946;
    wire _8947;
    wire _8948;
    wire _8949;
    wire _8950;
    wire _8951;
    wire _8952;
    wire _8953;
    wire _8954;
    wire _8955;
    wire _8956;
    wire _7795 = 1'b0;
    wire _7693;
    wire _7471 = 1'b0;
    wire _7469 = 1'b0;
    wire _7688 = 1'b1;
    wire _9014;
    wire _9015;
    wire _9016;
    wire _9017;
    wire _9018;
    wire _9019;
    wire _9020;
    wire _9021;
    wire _9022;
    wire _9023;
    wire _9024;
    wire _9025;
    wire _9026;
    wire _9027;
    wire _9028;
    wire _9029;
    wire _9030;
    wire _9031;
    wire _9032;
    wire _9033;
    wire _9034;
    wire _9035;
    wire _9036;
    wire _9037;
    wire _9038;
    wire _9039;
    wire _9040;
    wire _9041;
    wire _9042;
    wire _9043;
    wire _9044;
    wire [31:0] _7535 = 32'b00000000000000000000000000000000;
    wire [31:0] _7533 = 32'b00000000000000000000000000000000;
    wire _7571 = 1'b0;
    wire _7840;
    wire _8601;
    wire _8602;
    wire _8603;
    wire _8604;
    wire _8605;
    wire _8606;
    wire _8607;
    wire _8608;
    wire _8609;
    wire _8610;
    wire _7570;
    reg _7572;
    wire _7577 = 1'b0;
    wire _7842;
    wire _8581;
    wire _8582;
    wire _8583;
    wire _8584;
    wire _8585;
    wire _8586;
    wire _8587;
    wire _8588;
    wire _8589;
    wire _8590;
    wire _7576;
    reg _7578;
    wire _7580 = 1'b0;
    wire _7843;
    wire _8571;
    wire _8572;
    wire _8573;
    wire _8574;
    wire _8575;
    wire _8576;
    wire _8577;
    wire _8578;
    wire _8579;
    wire _8580;
    wire _7579;
    reg _7581;
    wire _7583 = 1'b0;
    wire _7844;
    wire _8561;
    wire _8562;
    wire _8563;
    wire _8564;
    wire _8565;
    wire _8566;
    wire _8567;
    wire _8568;
    wire _8569;
    wire _8570;
    wire _7582;
    reg _7584;
    wire _7586 = 1'b0;
    wire _7845;
    wire _8551;
    wire _8552;
    wire _8553;
    wire _8554;
    wire _8555;
    wire _8556;
    wire _8557;
    wire _8558;
    wire _8559;
    wire _8560;
    wire _7585;
    reg _7587;
    wire _7589 = 1'b0;
    wire _7846;
    wire _8541;
    wire _8542;
    wire _8543;
    wire _8544;
    wire _8545;
    wire _8546;
    wire _8547;
    wire _8548;
    wire _8549;
    wire _8550;
    wire _7588;
    reg _7590;
    wire _7592 = 1'b0;
    wire _7847;
    wire _8531;
    wire _8532;
    wire _8533;
    wire _8534;
    wire _8535;
    wire _8536;
    wire _8537;
    wire _8538;
    wire _8539;
    wire _8540;
    wire _7591;
    reg _7593;
    wire _7595 = 1'b0;
    wire _7848;
    wire _8521;
    wire _8522;
    wire _8523;
    wire _8524;
    wire _8525;
    wire _8526;
    wire _8527;
    wire _8528;
    wire _8529;
    wire _8530;
    wire _7594;
    reg _7596;
    wire _7598 = 1'b0;
    wire _7849;
    wire _8511;
    wire _8512;
    wire _8513;
    wire _8514;
    wire _8515;
    wire _8516;
    wire _8517;
    wire _8518;
    wire _8519;
    wire _8520;
    wire _7597;
    reg _7599;
    wire _7601 = 1'b0;
    wire _7850;
    wire _8501;
    wire _8502;
    wire _8503;
    wire _8504;
    wire _8505;
    wire _8506;
    wire _8507;
    wire _8508;
    wire _8509;
    wire _8510;
    wire _7600;
    reg _7602;
    wire _7604 = 1'b0;
    wire _7851;
    wire _8491;
    wire _8492;
    wire _8493;
    wire _8494;
    wire _8495;
    wire _8496;
    wire _8497;
    wire _8498;
    wire _8499;
    wire _8500;
    wire _7603;
    reg _7605;
    wire _7607 = 1'b0;
    wire _7852;
    wire _8481;
    wire _8482;
    wire _8483;
    wire _8484;
    wire _8485;
    wire _8486;
    wire _8487;
    wire _8488;
    wire _8489;
    wire _8490;
    wire _7606;
    reg _7608;
    wire _7610 = 1'b0;
    wire _7853;
    wire _8471;
    wire _8472;
    wire _8473;
    wire _8474;
    wire _8475;
    wire _8476;
    wire _8477;
    wire _8478;
    wire _8479;
    wire _8480;
    wire _7609;
    reg _7611;
    wire _7613 = 1'b0;
    wire _7854;
    wire _8461;
    wire _8462;
    wire _8463;
    wire _8464;
    wire _8465;
    wire _8466;
    wire _8467;
    wire _8468;
    wire _8469;
    wire _8470;
    wire _7612;
    reg _7614;
    wire _7616 = 1'b0;
    wire _7855;
    wire _8451;
    wire _8452;
    wire _8453;
    wire _8454;
    wire _8455;
    wire _8456;
    wire _8457;
    wire _8458;
    wire _8459;
    wire _8460;
    wire _7615;
    reg _7617;
    wire _7619 = 1'b0;
    wire _7856;
    wire _8441;
    wire _8442;
    wire _8443;
    wire _8444;
    wire _8445;
    wire _8446;
    wire _8447;
    wire _8448;
    wire _8449;
    wire _8450;
    wire _7618;
    reg _7620;
    wire _7622 = 1'b0;
    wire _7857;
    wire _8431;
    wire _8432;
    wire _8433;
    wire _8434;
    wire _8435;
    wire _8436;
    wire _8437;
    wire _8438;
    wire _8439;
    wire _8440;
    wire _7621;
    reg _7623;
    wire _7625 = 1'b0;
    wire _7858;
    wire _8421;
    wire _8422;
    wire _8423;
    wire _8424;
    wire _8425;
    wire _8426;
    wire _8427;
    wire _8428;
    wire _8429;
    wire _8430;
    wire _7624;
    reg _7626;
    wire _7628 = 1'b0;
    wire _7859;
    wire _8411;
    wire _8412;
    wire _8413;
    wire _8414;
    wire _8415;
    wire _8416;
    wire _8417;
    wire _8418;
    wire _8419;
    wire _8420;
    wire _7627;
    reg _7629;
    wire _7631 = 1'b0;
    wire _7860;
    wire _8401;
    wire _8402;
    wire _8403;
    wire _8404;
    wire _8405;
    wire _8406;
    wire _8407;
    wire _8408;
    wire _8409;
    wire _8410;
    wire _7630;
    reg _7632;
    wire _7634 = 1'b0;
    wire _7861;
    wire _8391;
    wire _8392;
    wire _8393;
    wire _8394;
    wire _8395;
    wire _8396;
    wire _8397;
    wire _8398;
    wire _8399;
    wire _8400;
    wire _7633;
    reg _7635;
    wire _7637 = 1'b0;
    wire _7862;
    wire _8381;
    wire _8382;
    wire _8383;
    wire _8384;
    wire _8385;
    wire _8386;
    wire _8387;
    wire _8388;
    wire _8389;
    wire _8390;
    wire _7636;
    reg _7638;
    wire _7640 = 1'b0;
    wire _7863;
    wire _8371;
    wire _8372;
    wire _8373;
    wire _8374;
    wire _8375;
    wire _8376;
    wire _8377;
    wire _8378;
    wire _8379;
    wire _8380;
    wire _7639;
    reg _7641;
    wire _7643 = 1'b0;
    wire _7864;
    wire _8361;
    wire _8362;
    wire _8363;
    wire _8364;
    wire _8365;
    wire _8366;
    wire _8367;
    wire _8368;
    wire _8369;
    wire _8370;
    wire _7642;
    reg _7644;
    wire _7646 = 1'b0;
    wire _7865;
    wire _8351;
    wire _8352;
    wire _8353;
    wire _8354;
    wire _8355;
    wire _8356;
    wire _8357;
    wire _8358;
    wire _8359;
    wire _8360;
    wire _7645;
    reg _7647;
    wire _7649 = 1'b0;
    wire _7866;
    wire _8341;
    wire _8342;
    wire _8343;
    wire _8344;
    wire _8345;
    wire _8346;
    wire _8347;
    wire _8348;
    wire _8349;
    wire _8350;
    wire _7648;
    reg _7650;
    wire _7652 = 1'b0;
    wire _7867;
    wire _8331;
    wire _8332;
    wire _8333;
    wire _8334;
    wire _8335;
    wire _8336;
    wire _8337;
    wire _8338;
    wire _8339;
    wire _8340;
    wire _7651;
    reg _7653;
    wire _7655 = 1'b0;
    wire _7868;
    wire _8321;
    wire _8322;
    wire _8323;
    wire _8324;
    wire _8325;
    wire _8326;
    wire _8327;
    wire _8328;
    wire _8329;
    wire _8330;
    wire _7654;
    reg _7656;
    wire _7658 = 1'b0;
    wire _7869;
    wire _8311;
    wire _8312;
    wire _8313;
    wire _8314;
    wire _8315;
    wire _8316;
    wire _8317;
    wire _8318;
    wire _8319;
    wire _8320;
    wire _7657;
    reg _7659;
    wire _7661 = 1'b0;
    wire _7870;
    wire _8301;
    wire _8302;
    wire _8303;
    wire _8304;
    wire _8305;
    wire _8306;
    wire _8307;
    wire _8308;
    wire _8309;
    wire _8310;
    wire _7660;
    reg _7662;
    wire _7664 = 1'b0;
    wire _7871;
    wire _8291;
    wire _8292;
    wire _8293;
    wire _8294;
    wire _8295;
    wire _8296;
    wire _8297;
    wire _8298;
    wire _8299;
    wire _8300;
    wire _7663;
    reg _7665;
    wire [31:0] _7666;
    wire [31:0] _7796;
    wire [31:0] _8660;
    wire [31:0] _8661;
    wire [31:0] _8662;
    wire [31:0] _8663;
    wire _8086 = 1'b1;
    wire [31:0] _8089 = 32'b00000000000000000000000000000000;
    wire [31:0] _8087 = 32'b00000000000000000000000000000001;
    wire [31:0] _8088;
    wire _8090;
    wire _8658;
    wire _8105;
    wire _8106;
    wire _8107;
    wire _8108;
    wire _8109;
    wire _8657;
    wire [31:0] _8091 = 32'b00000000000000000000000000000000;
    wire [31:0] _7672 = 32'b00000000000000000000000000000000;
    wire [31:0] _7670 = 32'b00000000000000000000000000000000;
    wire [31:0] _8269;
    wire [31:0] _8270;
    wire [31:0] _8271;
    wire [31:0] _8272;
    wire [31:0] _8273;
    wire [31:0] _8274;
    wire [31:0] _8275;
    wire [31:0] _8276;
    wire [31:0] _8084 = 32'b00000000000000000000000000000001;
    wire [31:0] _8085;
    wire [31:0] _8268;
    wire _8277;
    wire [31:0] _8278;
    wire [31:0] _7671;
    reg [31:0] _7673;
    wire _8092;
    wire _8093;
    wire _8094;
    wire _8095;
    wire _8659;
    wire _7537;
    wire _7916 = 1'b1;
    wire _7917;
    wire _7918;
    wire _7919;
    wire _7920;
    wire _8642;
    wire _8643;
    wire _8644;
    wire _8645;
    wire _7911 = 1'b1;
    wire _7912;
    wire _7913;
    wire _7914;
    wire _7915;
    wire _8646;
    wire _8647;
    wire _8648;
    wire _7931 = 1'b1;
    wire _7932;
    wire _7574 = 1'b0;
    wire [31:0] _37 = 32'b00000000000000000000000000000000;
    wire _7376;
    wire _7377;
    wire [31:0] _7379 = 32'b00000000000000000000000000000000;
    wire [31:0] _7378 = 32'b00000000000000000000000000000000;
    reg [31:0] _7380;
    wire _7371;
    wire _7372;
    wire [31:0] _7374 = 32'b00000000000000000000000000000000;
    wire [31:0] _7373 = 32'b00000000000000000000000000000000;
    reg [31:0] _7375;
    wire _7366;
    wire _7367;
    wire [31:0] _7369 = 32'b00000000000000000000000000000000;
    wire [31:0] _7368 = 32'b00000000000000000000000000000000;
    reg [31:0] _7370;
    wire _7361;
    wire _7362;
    wire [31:0] _7364 = 32'b00000000000000000000000000000000;
    wire [31:0] _7363 = 32'b00000000000000000000000000000000;
    reg [31:0] _7365;
    wire _7356;
    wire _7357;
    wire [31:0] _7359 = 32'b00000000000000000000000000000000;
    wire [31:0] _7358 = 32'b00000000000000000000000000000000;
    reg [31:0] _7360;
    wire _7351;
    wire _7352;
    wire [31:0] _7354 = 32'b00000000000000000000000000000000;
    wire [31:0] _7353 = 32'b00000000000000000000000000000000;
    reg [31:0] _7355;
    wire _7346;
    wire _7347;
    wire [31:0] _7349 = 32'b00000000000000000000000000000000;
    wire [31:0] _7348 = 32'b00000000000000000000000000000000;
    reg [31:0] _7350;
    wire _7341;
    wire _7342;
    wire [31:0] _7344 = 32'b00000000000000000000000000000000;
    wire [31:0] _7343 = 32'b00000000000000000000000000000000;
    reg [31:0] _7345;
    wire _7336;
    wire _7337;
    wire [31:0] _7339 = 32'b00000000000000000000000000000000;
    wire [31:0] _7338 = 32'b00000000000000000000000000000000;
    reg [31:0] _7340;
    wire _7331;
    wire _7332;
    wire [31:0] _7334 = 32'b00000000000000000000000000000000;
    wire [31:0] _7333 = 32'b00000000000000000000000000000000;
    reg [31:0] _7335;
    wire _7326;
    wire _7327;
    wire [31:0] _7329 = 32'b00000000000000000000000000000000;
    wire [31:0] _7328 = 32'b00000000000000000000000000000000;
    reg [31:0] _7330;
    wire _7321;
    wire _7322;
    wire [31:0] _7324 = 32'b00000000000000000000000000000000;
    wire [31:0] _7323 = 32'b00000000000000000000000000000000;
    reg [31:0] _7325;
    wire _7316;
    wire _7317;
    wire [31:0] _7319 = 32'b00000000000000000000000000000000;
    wire [31:0] _7318 = 32'b00000000000000000000000000000000;
    reg [31:0] _7320;
    wire _7311;
    wire _7312;
    wire [31:0] _7314 = 32'b00000000000000000000000000000000;
    wire [31:0] _7313 = 32'b00000000000000000000000000000000;
    reg [31:0] _7315;
    wire _7306;
    wire _7307;
    wire [31:0] _7309 = 32'b00000000000000000000000000000000;
    wire [31:0] _7308 = 32'b00000000000000000000000000000000;
    reg [31:0] _7310;
    wire _7301;
    wire _7302;
    wire [31:0] _7304 = 32'b00000000000000000000000000000000;
    wire [31:0] _7303 = 32'b00000000000000000000000000000000;
    reg [31:0] _7305;
    wire _7296;
    wire _7297;
    wire [31:0] _7299 = 32'b00000000000000000000000000000000;
    wire [31:0] _7298 = 32'b00000000000000000000000000000000;
    reg [31:0] _7300;
    wire _7291;
    wire _7292;
    wire [31:0] _7294 = 32'b00000000000000000000000000000000;
    wire [31:0] _7293 = 32'b00000000000000000000000000000000;
    reg [31:0] _7295;
    wire _7286;
    wire _7287;
    wire [31:0] _7289 = 32'b00000000000000000000000000000000;
    wire [31:0] _7288 = 32'b00000000000000000000000000000000;
    reg [31:0] _7290;
    wire _7281;
    wire _7282;
    wire [31:0] _7284 = 32'b00000000000000000000000000000000;
    wire [31:0] _7283 = 32'b00000000000000000000000000000000;
    reg [31:0] _7285;
    wire _7276;
    wire _7277;
    wire [31:0] _7279 = 32'b00000000000000000000000000000000;
    wire [31:0] _7278 = 32'b00000000000000000000000000000000;
    reg [31:0] _7280;
    wire _7271;
    wire _7272;
    wire [31:0] _7274 = 32'b00000000000000000000000000000000;
    wire [31:0] _7273 = 32'b00000000000000000000000000000000;
    reg [31:0] _7275;
    wire _7266;
    wire _7267;
    wire [31:0] _7269 = 32'b00000000000000000000000000000000;
    wire [31:0] _7268 = 32'b00000000000000000000000000000000;
    reg [31:0] _7270;
    wire _7261;
    wire _7262;
    wire [31:0] _7264 = 32'b00000000000000000000000000000000;
    wire [31:0] _7263 = 32'b00000000000000000000000000000000;
    reg [31:0] _7265;
    wire _7256;
    wire _7257;
    wire [31:0] _7259 = 32'b00000000000000000000000000000000;
    wire [31:0] _7258 = 32'b00000000000000000000000000000000;
    reg [31:0] _7260;
    wire _7251;
    wire _7252;
    wire [31:0] _7254 = 32'b00000000000000000000000000000000;
    wire [31:0] _7253 = 32'b00000000000000000000000000000000;
    reg [31:0] _7255;
    wire _7246;
    wire _7247;
    wire [31:0] _7249 = 32'b00000000000000000000000000000000;
    wire [31:0] _7248 = 32'b00000000000000000000000000000000;
    reg [31:0] _7250;
    wire _7241;
    wire _7242;
    wire [31:0] _7244 = 32'b00000000000000000000000000000000;
    wire [31:0] _7243 = 32'b00000000000000000000000000000000;
    reg [31:0] _7245;
    wire _7236;
    wire _7237;
    wire [31:0] _7239 = 32'b00000000000000000000000000000000;
    wire [31:0] _7238 = 32'b00000000000000000000000000000000;
    reg [31:0] _7240;
    wire _7231;
    wire _7232;
    wire [31:0] _7234 = 32'b00000000000000000000000000000000;
    wire [31:0] _7233 = 32'b00000000000000000000000000000000;
    reg [31:0] _7235;
    wire _7226;
    wire _7227;
    wire [31:0] _7229 = 32'b00000000000000000000000000000000;
    wire [31:0] _7228 = 32'b00000000000000000000000000000000;
    reg [31:0] _7230;
    wire _7221;
    wire _7222;
    wire [31:0] _7224 = 32'b00000000000000000000000000000000;
    wire [31:0] _7223 = 32'b00000000000000000000000000000000;
    reg [31:0] _7225;
    wire _7216;
    wire _7217;
    wire [31:0] _7219 = 32'b00000000000000000000000000000000;
    wire [31:0] _7218 = 32'b00000000000000000000000000000000;
    reg [31:0] _7220;
    wire _7211;
    wire _7212;
    wire [31:0] _7214 = 32'b00000000000000000000000000000000;
    wire [31:0] _7213 = 32'b00000000000000000000000000000000;
    reg [31:0] _7215;
    wire _6817;
    wire _6820;
    wire _6828;
    wire _6848;
    wire _6896;
    wire _7008;
    wire _6818;
    wire _6819;
    wire _6827;
    wire _6847;
    wire _6895;
    wire _7007;
    wire _6821;
    wire _6823;
    wire _6826;
    wire _6846;
    wire _6894;
    wire _7006;
    wire _6822;
    wire _6824;
    wire _6825;
    wire _6845;
    wire _6893;
    wire _7005;
    wire _6829;
    wire _6832;
    wire _6839;
    wire _6844;
    wire _6892;
    wire _7004;
    wire _6830;
    wire _6831;
    wire _6838;
    wire _6843;
    wire _6891;
    wire _7003;
    wire _6833;
    wire _6835;
    wire _6837;
    wire _6842;
    wire _6890;
    wire _7002;
    wire _6834;
    wire _6836;
    wire _6840;
    wire _6841;
    wire _6889;
    wire _7001;
    wire _6849;
    wire _6852;
    wire _6860;
    wire _6879;
    wire _6888;
    wire _7000;
    wire _6850;
    wire _6851;
    wire _6859;
    wire _6878;
    wire _6887;
    wire _6999;
    wire _6853;
    wire _6855;
    wire _6858;
    wire _6877;
    wire _6886;
    wire _6998;
    wire _6854;
    wire _6856;
    wire _6857;
    wire _6876;
    wire _6885;
    wire _6997;
    wire _6861;
    wire _6864;
    wire _6871;
    wire _6875;
    wire _6884;
    wire _6996;
    wire _6862;
    wire _6863;
    wire _6870;
    wire _6874;
    wire _6883;
    wire _6995;
    wire _6865;
    wire _6867;
    wire _6869;
    wire _6873;
    wire _6882;
    wire _6994;
    wire _6866;
    wire _6868;
    wire _6872;
    wire _6880;
    wire _6881;
    wire _6993;
    wire _6897;
    wire _6900;
    wire _6908;
    wire _6928;
    wire _6975;
    wire _6992;
    wire _6898;
    wire _6899;
    wire _6907;
    wire _6927;
    wire _6974;
    wire _6991;
    wire _6901;
    wire _6903;
    wire _6906;
    wire _6926;
    wire _6973;
    wire _6990;
    wire _6902;
    wire _6904;
    wire _6905;
    wire _6925;
    wire _6972;
    wire _6989;
    wire _6909;
    wire _6912;
    wire _6919;
    wire _6924;
    wire _6971;
    wire _6988;
    wire _6910;
    wire _6911;
    wire _6918;
    wire _6923;
    wire _6970;
    wire _6987;
    wire _6913;
    wire _6915;
    wire _6917;
    wire _6922;
    wire _6969;
    wire _6986;
    wire _6914;
    wire _6916;
    wire _6920;
    wire _6921;
    wire _6968;
    wire _6985;
    wire _6929;
    wire _6932;
    wire _6940;
    wire _6959;
    wire _6967;
    wire _6984;
    wire _6930;
    wire _6931;
    wire _6939;
    wire _6958;
    wire _6966;
    wire _6983;
    wire _6933;
    wire _6935;
    wire _6938;
    wire _6957;
    wire _6965;
    wire _6982;
    wire _6934;
    wire _6936;
    wire _6937;
    wire _6956;
    wire _6964;
    wire _6981;
    wire _6941;
    wire _6944;
    wire _6951;
    wire _6955;
    wire _6963;
    wire _6980;
    wire _6942;
    wire _6943;
    wire _6950;
    wire _6954;
    wire _6962;
    wire _6979;
    wire _6945;
    wire _6947;
    wire _6949;
    wire _6953;
    wire _6961;
    wire _6978;
    wire _6946;
    wire _6948;
    wire _6952;
    wire _6960;
    wire _6976;
    wire _6977;
    wire _7009;
    wire _7012;
    wire _7020;
    wire _7040;
    wire _7088;
    wire _7199;
    wire _7010;
    wire _7011;
    wire _7019;
    wire _7039;
    wire _7087;
    wire _7198;
    wire _7013;
    wire _7015;
    wire _7018;
    wire _7038;
    wire _7086;
    wire _7197;
    wire _7014;
    wire _7016;
    wire _7017;
    wire _7037;
    wire _7085;
    wire _7196;
    wire _7021;
    wire _7024;
    wire _7031;
    wire _7036;
    wire _7084;
    wire _7195;
    wire _7022;
    wire _7023;
    wire _7030;
    wire _7035;
    wire _7083;
    wire _7194;
    wire _7025;
    wire _7027;
    wire _7029;
    wire _7034;
    wire _7082;
    wire _7193;
    wire _7026;
    wire _7028;
    wire _7032;
    wire _7033;
    wire _7081;
    wire _7192;
    wire _7041;
    wire _7044;
    wire _7052;
    wire _7071;
    wire _7080;
    wire _7191;
    wire _7042;
    wire _7043;
    wire _7051;
    wire _7070;
    wire _7079;
    wire _7190;
    wire _7045;
    wire _7047;
    wire _7050;
    wire _7069;
    wire _7078;
    wire _7189;
    wire _7046;
    wire _7048;
    wire _7049;
    wire _7068;
    wire _7077;
    wire _7188;
    wire _7053;
    wire _7056;
    wire _7063;
    wire _7067;
    wire _7076;
    wire _7187;
    wire _7054;
    wire _7055;
    wire _7062;
    wire _7066;
    wire _7075;
    wire _7186;
    wire _7057;
    wire _7059;
    wire _7061;
    wire _7065;
    wire _7074;
    wire _7185;
    wire _7058;
    wire _7060;
    wire _7064;
    wire _7072;
    wire _7073;
    wire _7184;
    wire _7089;
    wire _7092;
    wire _7100;
    wire _7120;
    wire _7167;
    wire _7183;
    wire _7090;
    wire _7091;
    wire _7099;
    wire _7119;
    wire _7166;
    wire _7182;
    wire _7093;
    wire _7095;
    wire _7098;
    wire _7118;
    wire _7165;
    wire _7181;
    wire _7094;
    wire _7096;
    wire _7097;
    wire _7117;
    wire _7164;
    wire _7180;
    wire _7101;
    wire _7104;
    wire _7111;
    wire _7116;
    wire _7163;
    wire _7179;
    wire _7102;
    wire _7103;
    wire _7110;
    wire _7115;
    wire _7162;
    wire _7178;
    wire _7105;
    wire _7107;
    wire _7109;
    wire _7114;
    wire _7161;
    wire _7177;
    wire _7106;
    wire _7108;
    wire _7112;
    wire _7113;
    wire _7160;
    wire _7176;
    wire _7121;
    wire _7124;
    wire _7132;
    wire _7151;
    wire _7159;
    wire _7175;
    wire _7122;
    wire _7123;
    wire _7131;
    wire _7150;
    wire _7158;
    wire _7174;
    wire _7125;
    wire _7127;
    wire _7130;
    wire _7149;
    wire _7157;
    wire _7173;
    wire _7126;
    wire _7128;
    wire _7129;
    wire _7148;
    wire _7156;
    wire _7172;
    wire _7133;
    wire _7136;
    wire _7143;
    wire _7147;
    wire _7155;
    wire _7171;
    wire _7134;
    wire _7135;
    wire _7142;
    wire _7146;
    wire _7154;
    wire _7170;
    wire _7137;
    wire _7139;
    wire _7141;
    wire _7145;
    wire _7153;
    wire _7169;
    wire _6811;
    wire _6812;
    wire _7138;
    wire _6813;
    wire _7140;
    wire _6814;
    wire _7144;
    wire _6815;
    wire _7152;
    wire [5:0] _6806 = 6'b000000;
    wire [5:0] _6804 = 6'b000000;
    wire _7700;
    wire [4:0] _7703 = 5'b00000;
    wire [5:0] _7705;
    wire [5:0] _7706 = 6'b100000;
    wire [5:0] _7707;
    wire [5:0] _7698 = 6'b000100;
    wire [5:0] _7697 = 6'b000011;
    wire _7699;
    wire [5:0] _9113;
    wire [5:0] _9114;
    wire [4:0] _6557 = 5'b00000;
    wire [4:0] _6556 = 5'b00000;
    wire [4:0] _6555;
    reg [4:0] _6558;
    wire [5:0] _6559;
    wire [5:0] _5642;
    wire [5:0] _9115;
    wire [5:0] _7882 = 6'b100000;
    wire [5:0] _7883;
    wire [5:0] _9116;
    wire [5:0] _9117;
    wire [5:0] _9118;
    wire [5:0] _9119;
    wire [5:0] _9120;
    wire [5:0] _7947 = 6'b000000;
    wire [5:0] _9121;
    wire _9122;
    wire [5:0] _9123;
    wire _9124;
    wire [5:0] _9125;
    wire _9126;
    wire [5:0] _9127;
    wire [5:0] _6805;
    reg [5:0] _6807;
    wire _6816;
    wire _7168;
    wire [63:0] _7200;
    wire _7206;
    wire _9093;
    wire _9094;
    wire _9095;
    wire _9096;
    wire _7801;
    wire _7802;
    wire _9097;
    wire [1:0] _7527 = 2'b00;
    wire [1:0] _7525 = 2'b00;
    wire [1:0] _7713 = 2'b01;
    wire [1:0] _7709 = 2'b10;
    wire [1:0] _7708 = 2'b00;
    wire [1:0] _7710 = 2'b01;
    wire _7711;
    wire [1:0] _7712;
    wire [1:0] _7714 = 2'b00;
    wire _7715;
    wire [1:0] _7716;
    wire [1:0] _8679;
    wire _8680;
    wire [1:0] _8681;
    wire [1:0] _7526;
    reg [1:0] _7528;
    wire _7805;
    wire _7806;
    wire _9098;
    wire _9099;
    wire _9100;
    wire _9101;
    wire _9102;
    wire _6810;
    wire _7207;
    wire [31:0] _7209 = 32'b00000000000000000000000000000000;
    wire [31:0] _7208 = 32'b00000000000000000000000000000000;
    reg [31:0] _7210;
    reg [31:0] _7382;
    wire [31:0] _7816 = 32'b00000000000000000000000000000000;
    wire [5:0] _7817 = 6'b000000;
    wire [5:0] _6553 = 6'b000000;
    wire [5:0] _6552 = 6'b000000;
    wire [5:0] _6469 = 6'b100000;
    wire [4:0] _6466;
    wire [5:0] _6467;
    wire [4:0] _6464;
    wire [5:0] cx;
    wire [6:0] _6448 = 7'b0000000;
    wire [6:0] _6447;
    wire _6449;
    wire [6:0] _6451 = 7'b0001011;
    wire [6:0] _6450;
    wire _6452;
    wire _6453;
    wire _6454;
    wire c0;
    wire [5:0] _6468;
    wire [6:0] _6457 = 7'b0000010;
    wire [6:0] _6456;
    wire _6458;
    wire [6:0] _6460 = 7'b0001011;
    wire [6:0] _6459;
    wire _6461;
    wire _6462;
    wire c1;
    wire [5:0] _6470;
    reg [5:0] _6554;
    wire [5:0] _5641;
    wire _7818;
    wire _7819;
    wire [31:0] _7820;
    wire [31:0] _7839;
    wire _7841;
    wire _8591;
    wire _8592;
    wire _8593;
    wire _8594;
    wire _8595;
    wire _8596;
    wire _8597;
    wire _8598;
    wire _8599;
    wire _8600;
    wire _7573;
    reg _7575;
    wire _7933;
    wire _7934;
    wire _7935;
    wire _8649;
    wire _7463 = 1'b0;
    wire _7461 = 1'b0;
    wire [3:0] _8098 = 4'b0000;
    wire [3:0] _7467 = 4'b0000;
    wire [3:0] _7465 = 4'b0000;
    wire [3:0] _8101 = 4'b0001;
    wire [3:0] _8102;
    wire _9082;
    wire _9083;
    wire _9084;
    wire _9085;
    wire _9086;
    wire _9087;
    wire _9088;
    wire [3:0] _9089;
    wire [3:0] _8100 = 4'b1111;
    wire _5830;
    wire _5831;
    wire _5832;
    wire _5635;
    wire _8103;
    wire _8104;
    wire [3:0] _9090;
    wire [3:0] _9091;
    wire [3:0] _7466;
    reg [3:0] _7468;
    wire _8099;
    wire _9092;
    wire _7462;
    reg _7464;
    wire _8650;
    wire _8651;
    wire _8652;
    wire _8110;
    wire _8111;
    wire _8112;
    wire _8113;
    wire _8114;
    wire _8641;
    wire _8653;
    wire _8654;
    wire _8655;
    wire _8656;
    wire _7538;
    wire _8115;
    wire _8116;
    wire _8117;
    wire _8118;
    wire _8119;
    wire _8640;
    wire _7539;
    wire _8120;
    wire _8121;
    wire _8122;
    wire _8123;
    wire _8124;
    wire _8639;
    wire _7540;
    wire _8125;
    wire _8126;
    wire _8127;
    wire _8128;
    wire _8129;
    wire _8638;
    wire _7541;
    wire _8130;
    wire _8131;
    wire _8132;
    wire _8133;
    wire _8134;
    wire _8637;
    wire _7542;
    wire _8135;
    wire _8136;
    wire _8137;
    wire _8138;
    wire _8139;
    wire _8636;
    wire _7543;
    wire _8140;
    wire _8141;
    wire _8142;
    wire _8143;
    wire _8144;
    wire _8635;
    wire _7544;
    wire _8145;
    wire _8146;
    wire _8147;
    wire _8148;
    wire _8149;
    wire _8634;
    wire _7545;
    wire _8150;
    wire _8151;
    wire _8152;
    wire _8153;
    wire _8154;
    wire _8633;
    wire _7546;
    wire _8155;
    wire _8156;
    wire _8157;
    wire _8158;
    wire _8159;
    wire _8632;
    wire _7547;
    wire _8160;
    wire _8161;
    wire _8162;
    wire _8163;
    wire _8164;
    wire _8631;
    wire _7548;
    wire _8165;
    wire _8166;
    wire _8167;
    wire _8168;
    wire _8169;
    wire _8630;
    wire _7549;
    wire _8170;
    wire _8171;
    wire _8172;
    wire _8173;
    wire _8174;
    wire _8629;
    wire _7550;
    wire _8175;
    wire _8176;
    wire _8177;
    wire _8178;
    wire _8179;
    wire _8628;
    wire _7551;
    wire _8180;
    wire _8181;
    wire _8182;
    wire _8183;
    wire _8184;
    wire _8627;
    wire _7552;
    wire _8185;
    wire _8186;
    wire _8187;
    wire _8188;
    wire _8189;
    wire _8626;
    wire _7553;
    wire _8190;
    wire _8191;
    wire _8192;
    wire _8193;
    wire _8194;
    wire _8625;
    wire _7554;
    wire _8195;
    wire _8196;
    wire _8197;
    wire _8198;
    wire _8199;
    wire _8624;
    wire _7555;
    wire _8200;
    wire _8201;
    wire _8202;
    wire _8203;
    wire _8204;
    wire _8623;
    wire _7556;
    wire _8205;
    wire _8206;
    wire _8207;
    wire _8208;
    wire _8209;
    wire _8622;
    wire _7557;
    wire _8210;
    wire _8211;
    wire _8212;
    wire _8213;
    wire _8214;
    wire _8621;
    wire _7558;
    wire _8215;
    wire _8216;
    wire _8217;
    wire _8218;
    wire _8219;
    wire _8620;
    wire _7559;
    wire _8220;
    wire _8221;
    wire _8222;
    wire _8223;
    wire _8224;
    wire _8619;
    wire _7560;
    wire _8225;
    wire _8226;
    wire _8227;
    wire _8228;
    wire _8229;
    wire _8618;
    wire _7561;
    wire _8230;
    wire _8231;
    wire _8232;
    wire _8233;
    wire _8234;
    wire _8617;
    wire _7562;
    wire _8235;
    wire _8236;
    wire _8237;
    wire _8238;
    wire _8239;
    wire _8616;
    wire _7563;
    wire _8240;
    wire _8241;
    wire _8242;
    wire _8243;
    wire _8244;
    wire _8615;
    wire _7564;
    wire _8245;
    wire _8246;
    wire _8247;
    wire _8248;
    wire _8249;
    wire _8614;
    wire _7565;
    wire _8250;
    wire _8251;
    wire _8252;
    wire _8253;
    wire _8254;
    wire _8613;
    wire _7566;
    wire _8255;
    wire _8256;
    wire _8257;
    wire _8258;
    wire _8259;
    wire _8612;
    wire _7567;
    wire _8260;
    wire [31:0] _38 = 32'b11111111111111111111111111111111;
    wire _8261;
    wire _8262;
    wire _8263;
    wire _8264;
    wire _8611;
    wire _7568;
    wire [31:0] _7569;
    wire _8664;
    wire [31:0] _8665;
    wire [31:0] _7534;
    reg [31:0] _7536;
    wire _9045;
    wire _9046;
    wire _9047;
    wire _9048;
    wire _9049;
    wire _9050;
    wire _9051;
    wire _9052;
    wire _9053;
    wire _9054;
    wire _9055;
    wire _9056;
    wire _9057;
    wire _9058;
    wire _9059;
    wire _9060;
    wire _9061;
    wire _9062;
    wire _9063;
    wire _9064;
    wire _9065;
    wire _9066;
    wire _9067;
    wire _9068;
    wire _9069;
    wire _9070;
    wire _9071;
    wire _9072;
    wire _9073;
    wire _9074;
    wire _9075;
    wire _9076;
    wire _9077;
    wire _9078;
    wire _9079;
    wire _8081 = 1'b0;
    wire _9080;
    wire _9081;
    wire _7470;
    reg _7472;
    wire _7694;
    wire _7695;
    wire _7696;
    wire _8957;
    wire _8958;
    wire _8959;
    wire _8960;
    wire _8961;
    wire _7895 = 1'b1;
    wire _7887 = 1'b1;
    wire _7881 = 1'b1;
    wire _7875 = 1'b1;
    wire _7872 = 1'b1;
    wire _7835 = 1'b1;
    wire _7836;
    wire _7837;
    wire _7838;
    wire _8962;
    wire _7873;
    wire _7874;
    wire _8963;
    wire _8964;
    wire _8965;
    wire _8966;
    wire _8967;
    wire _8968;
    wire _8969;
    wire _5820 = 1'b0;
    reg _5821;
    wire _5836;
    wire _5837;
    wire _5637;
    wire _5822 = 1'b0;
    wire _5768 = 1'b0;
    wire _5811;
    wire _5765 = 1'b0;
    wire _5720 = 1'b0;
    reg _5721;
    wire _5722;
    wire _5718 = 1'b0;
    wire _5692 = 1'b0;
    wire [2:0] _5689 = 3'b000;
    wire [2:0] _5688;
    wire _5690;
    wire _5691;
    reg _5693;
    wire _5712;
    wire _5713;
    wire _5714;
    reg _5719;
    wire _5723;
    wire _5773;
    wire [6:0] _5762 = 7'b0000000;
    wire [6:0] _5760 = 7'b0000000;
    wire [6:0] _5775 = 7'b0111110;
    wire [6:0] _5774 = 7'b0011110;
    wire _5710 = 1'b0;
    wire [2:0] _5707 = 3'b011;
    wire [2:0] _5706;
    wire _5708;
    wire _5709;
    reg _5711;
    wire _5704 = 1'b0;
    wire [2:0] _5701 = 3'b010;
    wire [2:0] _5700;
    wire _5702;
    wire _5703;
    reg _5705;
    wire _5698 = 1'b0;
    wire [2:0] _5695 = 3'b001;
    wire [2:0] _5694;
    wire _5696;
    wire [6:0] _5680 = 7'b0000001;
    wire [6:0] _5679;
    wire _5681;
    wire [6:0] _5683 = 7'b0110011;
    wire [31:0] _6561 = 32'b00000000000000000000000000000000;
    wire [31:0] _6560 = 32'b00000000000000000000000000000000;
    reg [31:0] _6562;
    wire [31:0] _5643;
    wire [6:0] _5682;
    wire _5684;
    wire _6766 = 1'b0;
    wire _6764 = 1'b0;
    wire _7921 = 1'b0;
    wire _7924 = 1'b1;
    wire _9295;
    wire _9296;
    wire _9297;
    wire _9298;
    wire _7936 = 1'b0;
    wire _7938 = 1'b1;
    wire _9299;
    wire _9300;
    wire _9301;
    wire _9302;
    wire _9303;
    wire _9304;
    wire _6765;
    reg _6767;
    wire _5665;
    wire _5685;
    wire _5686;
    wire _5687;
    wire _5697;
    reg _5699;
    wire _5715;
    wire _5716;
    wire [6:0] _5776;
    wire [6:0] _5771 = 7'b0000001;
    wire [6:0] _5772;
    wire [6:0] _5815;
    wire [6:0] _5761;
    reg [6:0] _5763;
    wire _5770;
    wire _5813;
    wire _5814;
    wire _5764;
    reg _5766;
    wire _5812;
    wire _5767;
    reg _5769;
    reg _5823;
    wire _5833;
    wire _5834;
    wire _5835;
    wire _5634;
    wire _8970;
    wire _7939;
    wire _7940;
    wire _8971;
    wire _7943 = 1'b1;
    wire _8972;
    wire _8006 = 1'b1;
    wire _8073 = 1'b1;
    wire _8973;
    wire _8974;
    wire _8975;
    wire _8976;
    wire _8977;
    wire _8978;
    wire _8979;
    wire _8980;
    wire _8981;
    wire _8982;
    wire _8983;
    wire _8984;
    wire _7490;
    reg _7492;
    wire _8667;
    wire _8668;
    wire _7877 = 1'b0;
    wire _8669;
    wire _8670;
    wire _8671;
    wire _8672;
    wire _8673;
    wire _8674;
    wire _8675;
    wire _8676;
    wire _8677;
    wire _8678;
    wire _7530;
    reg _7532;
    wire _7785;
    wire _7786;
    wire _7787;
    wire _7788;
    wire _7789;
    wire _8993;
    wire _7876 = 1'b1;
    wire _7879;
    wire _7880;
    wire _8994;
    wire _7884;
    wire _7885;
    wire _7886;
    wire _8995;
    wire _7888;
    wire _7889;
    wire _7890;
    wire _8996;
    wire _7894;
    wire _8997;
    wire _7910;
    wire _8998;
    wire _7925;
    wire _8999;
    wire _7944;
    wire _9000;
    wire _9001;
    wire _9002;
    wire _9003;
    wire _9004;
    wire _9005;
    wire _9006;
    wire _7482;
    reg _7484;
    wire [31:0] _9110;
    wire [31:0] _6808 = 32'b00000000000000000000000000000000;
    wire _9111;
    wire [31:0] _9112;
    wire [31:0] _6809;
    reg [31:0] _7205;
    reg [31:0] _7381;
    wire [31:0] _7821 = 32'b00000000000000000000000000000000;
    wire [5:0] _7822 = 6'b000000;
    wire [4:0] _6549 = 5'b00000;
    wire [4:0] _6548 = 5'b00000;
    wire [4:0] _6547;
    reg [4:0] _6550;
    wire [5:0] _6551;
    wire [5:0] _5640;
    wire _7823;
    wire _7824;
    wire [31:0] _7825;
    wire [4:0] _7941;
    wire [4:0] _7974 = 5'b00100;
    wire [4:0] _7975;
    wire [4:0] _7950 = 5'b00001;
    wire [4:0] _7951;
    wire [4:0] _8001 = 5'b00100;
    wire _8002;
    wire _8003;
    wire [4:0] _8696;
    wire [4:0] _8697;
    wire [4:0] _8266 = 5'b00000;
    wire _8698;
    wire [4:0] _8699;
    wire _8700;
    wire [4:0] _8701;
    wire _8702;
    wire [4:0] _8703;
    wire [4:0] _7522;
    reg [4:0] _7524;
    wire _8005;
    wire [31:0] _9138;
    wire [31:0] _8012;
    wire [31:0] _9139;
    wire [31:0] _9140;
    wire _6754 = 1'b0;
    wire _6752 = 1'b0;
    wire _8007 = 1'b1;
    wire _9317;
    wire _9318;
    wire _8026 = 1'b1;
    wire _9319;
    wire _9320;
    wire _8082 = 1'b0;
    wire _9321;
    wire _9322;
    wire _9323;
    wire _9324;
    wire _6753;
    reg _6755;
    wire _5662;
    wire _5842;
    wire _5843;
    wire [31:0] _6545 = 32'b00000000000000000000000000000000;
    wire [31:0] _6544 = 32'b00000000000000000000000000000000;
    wire _5841;
    wire [31:0] _6488 = 32'b00000000000000000000000000000000;
    wire [31:0] _6487 = 32'b00000000000000000000000000000000;
    wire _6485;
    wire [9:0] _6482;
    wire _6483;
    wire [7:0] _6484;
    wire [2:0] _6475;
    wire [19:0] _6471;
    wire [20:0] _6472;
    wire _6473;
    wire [1:0] _6474;
    wire [3:0] _6476;
    wire [7:0] _6477;
    wire [10:0] _6478;
    wire [31:0] _6480;
    wire [11:0] _6481;
    wire [31:0] _6486;
    reg [31:0] _6489;
    wire [11:0] _6532 = 12'b000000000000;
    wire [19:0] _6533;
    wire [31:0] _6534;
    wire [11:0] _6518;
    wire _6519;
    wire [1:0] _6520;
    wire [3:0] _6521;
    wire [7:0] _6522;
    wire [15:0] _6523;
    wire [19:0] _6524;
    wire [31:0] _6526;
    wire [2:0] _6510;
    wire [3:0] _6506;
    wire [5:0] _6505;
    wire _6504;
    wire _6503;
    wire [12:0] _6507;
    wire _6508;
    wire [1:0] _6509;
    wire [3:0] _6511;
    wire [7:0] _6512;
    wire [15:0] _6513;
    wire [18:0] _6514;
    wire [31:0] _6516;
    wire [4:0] _6492;
    wire [6:0] _6491;
    wire [11:0] _6493;
    wire _6494;
    wire [1:0] _6495;
    wire [3:0] _6496;
    wire [7:0] _6497;
    wire [15:0] _6498;
    wire [19:0] _6499;
    wire [31:0] _6501;
    wire [31:0] _6490 = 32'b00000000000000000000000000000000;
    wire _6502;
    wire [31:0] _6539;
    wire _6517;
    wire [31:0] _6540;
    wire _6528;
    wire _6527;
    wire _6529;
    wire _6530;
    wire _6531;
    wire [31:0] _6541;
    wire _6536;
    wire _6535;
    wire _6537;
    wire [31:0] _6542;
    wire _6538;
    wire [31:0] _6543;
    reg [31:0] _6546;
    wire [31:0] _5639;
    wire [31:0] _8052;
    wire [31:0] _9141;
    wire [31:0] _9142;
    wire _9143;
    wire [31:0] _9144;
    wire _9145;
    wire [31:0] _9146;
    wire _9147;
    wire [31:0] _9148;
    wire _9149;
    wire [31:0] _9150;
    wire [31:0] _6797;
    reg [31:0] _6799;
    wire _7383;
    wire _7394;
    wire _7414;
    wire _7397;
    wire _7408;
    wire _7417;
    wire _7411;
    wire [47:0] _5645;
    wire _7413;
    wire _7419;
    wire _7421;
    wire _7422;
    wire _9305;
    wire _9306;
    wire _8008 = 1'b1;
    wire _8009;
    wire _8010;
    wire _9307;
    wire _9308;
    wire _8027 = 1'b1;
    wire _8049;
    wire _8050;
    wire _9309;
    wire _9310;
    wire _8083;
    wire _9311;
    wire _9312;
    wire _9313;
    wire _9314;
    wire _9315;
    wire _9316;
    wire _6761;
    reg _6763;
    wire _5664;
    wire _5846;
    wire _6239 = 1'b0;
    wire [2:0] _6236 = 3'b000;
    wire [31:0] _5652;
    wire [2:0] _6235;
    wire _6237;
    wire _5870 = 1'b0;
    wire [6:0] _5868 = 7'b1100011;
    wire [6:0] _5867;
    wire _5869;
    reg is_beq_bne_blt_bge_bltu_bgeu;
    wire _6238;
    reg instr_beq;
    wire _6249 = 1'b0;
    wire [6:0] _6242 = 7'b0000100;
    wire [6:0] _6241;
    wire _6243;
    wire [6:0] _6245 = 7'b0001011;
    wire [6:0] _6244;
    wire _6246;
    wire _6247;
    wire _6248;
    reg instr_waitirq;
    wire _6259 = 1'b0;
    wire [6:0] _6252 = 7'b0000010;
    wire [6:0] _6251;
    wire _6253;
    wire [6:0] _6255 = 7'b0001011;
    wire [6:0] _6254;
    wire _6256;
    wire _6257;
    wire _6258;
    reg instr_retirq;
    wire _5865 = 1'b0;
    wire [6:0] _5863 = 7'b1100111;
    wire [6:0] _5862;
    wire _5864;
    reg instr_jalr;
    wire _5860 = 1'b0;
    wire [6:0] _5858 = 7'b1101111;
    wire [6:0] _5857;
    wire _5859;
    reg instr_jal;
    wire _5855 = 1'b0;
    wire [6:0] _5853 = 7'b0010111;
    wire [6:0] _5852;
    wire _5854;
    reg instr_auipc;
    wire _5844;
    wire _5850 = 1'b0;
    wire [6:0] _5848 = 7'b0110111;
    wire _6599;
    wire [31:0] _6601 = 32'b00000000000000000000000000000000;
    wire [31:0] _6600 = 32'b00000000000000000000000000000000;
    reg [31:0] _6602;
    wire _6576 = 1'b0;
    wire _6778 = 1'b0;
    wire _6776 = 1'b0;
    wire _8075 = 1'b1;
    wire _8078 = 1'b0;
    wire _9276;
    wire _8051 = 1'b1;
    wire _8070;
    wire _8283;
    wire _8284;
    wire _8285;
    wire _8286;
    wire _7668;
    wire _9277;
    wire _6777;
    reg _6779;
    wire _5668;
    wire _5666;
    wire _6695;
    wire _6696;
    wire _6708;
    wire vdd = 1'b1;
    wire _6782 = 1'b0;
    wire _6780 = 1'b0;
    wire _8074 = 1'b1;
    wire _8077 = 1'b0;
    wire _9274;
    wire _8011 = 1'b1;
    wire _8023;
    wire _8287;
    wire _8024;
    wire _8025;
    wire _8288;
    wire _8289;
    wire _8290;
    wire _7667;
    wire _9275;
    wire _6781;
    reg _6783;
    wire _5669;
    wire _6709;
    wire _6710;
    wire _6711;
    wire _6712;
    wire _6713;
    wire _6714;
    wire _6715;
    wire _6716;
    wire _6717;
    wire _6575;
    reg _6577;
    wire _6603;
    wire _6604;
    wire [31:0] _6605;
    wire [31:0] _6598;
    wire [31:0] _5653;
    wire [6:0] _5847;
    wire _5849;
    reg instr_lui;
    wire _6261;
    wire _6262;
    wire _6263;
    wire _6264;
    wire _6265;
    wire _6266;
    wire _6267;
    wire _6268;
    wire _6269;
    wire _6270;
    wire _6271;
    wire _6272;
    wire _6273;
    wire _6274;
    wire _6275;
    wire _6276;
    wire _6277;
    wire _6278;
    wire _6279;
    wire _6280;
    wire _6281;
    wire _6282;
    wire _6283;
    wire _6284;
    wire _6285;
    wire _6286;
    wire _6287;
    wire _6288;
    wire _6289;
    wire _6290;
    wire _6291;
    wire _6292;
    wire _6293;
    wire _6294;
    wire _6295;
    wire _6296;
    wire _6297;
    wire _6298;
    wire _6299;
    wire _6300;
    wire _6301;
    wire _6302;
    wire _6303;
    wire _6304;
    wire _6305;
    wire _6306;
    wire instr_trap;
    wire [47:0] _6308;
    wire _6309;
    wire _6313;
    wire _6314;
    wire is_rdcycle_rdcycleh_rdinstr_rdinstrh;
    wire [14:0] _6446;
    wire [14:0] _5644;
    wire _7948;
    wire _8280;
    wire gnd = 1'b0;
    wire _8281;
    wire _8282;
    wire _7669;
    wire _9273;
    wire _6785;
    reg _6787;
    wire _5670;
    wire [1:0] _6723;
    wire [1:0] _6564 = 2'b11;
    wire _6724;
    wire [1:0] _6725;
    wire [1:0] _6565 = 2'b10;
    wire _6726;
    wire [1:0] _6727;
    wire [1:0] _6566 = 2'b01;
    wire _6728;
    wire [1:0] _6729;
    wire _6730;
    wire [1:0] _6731;
    wire [1:0] _6568;
    reg [1:0] _6570;
    wire [1:0] _6567 = 2'b00;
    wire _6573;
    wire _6574;
    wire _6584;
    wire _6585;
    wire _6586;
    wire _5659;
    wire _9294;
    wire _6769;
    reg _6771;
    wire _8071;
    wire _8072;
    wire [2:0] _9375;
    wire [2:0] _6733 = 3'b111;
    wire _9376;
    wire [2:0] _9377;
    wire [2:0] _6734 = 3'b110;
    wire _9378;
    wire [2:0] _9379;
    wire [2:0] _6735 = 3'b101;
    wire _9380;
    wire [2:0] _9381;
    wire [2:0] _6736 = 3'b100;
    wire _9382;
    wire [2:0] _9383;
    wire [2:0] _6737 = 3'b011;
    wire _9384;
    wire [2:0] _9385;
    wire [2:0] _6738 = 3'b010;
    wire _9386;
    wire [2:0] _9387;
    wire [2:0] _6740 = 3'b000;
    wire _9388;
    wire [2:0] _9389;
    wire [2:0] _6741;
    reg [2:0] _6743;
    wire _9169;
    wire _9170;
    wire _6789;
    reg _6791;
    wire _5671;

    /* logic */
    assign _7799 = ~ _7666;
    assign _7800 = _7536 & _7799;
    assign _9325 = _7802 ? _7800 : _6751;
    assign _9326 = _7806 ? _6751 : _9325;
    assign _9327 = _7492 ? _6751 : _9326;
    assign _9328 = _7484 ? _6751 : _9327;
    assign _9329 = _7880 ? _7878 : _6751;
    assign _9330 = _7886 ? _6751 : _9329;
    assign _9331 = _7890 ? _6751 : _9330;
    assign _9332 = _7894 ? _6751 : _9331;
    assign _9333 = _7910 ? _6751 : _9332;
    assign _9334 = _7925 ? _6751 : _9333;
    assign _9335 = _6743 == _6738;
    assign _9336 = _9335 ? _9334 : _6751;
    assign _9337 = _6743 == _6740;
    assign _9338 = _9337 ? _9328 : _9336;
    assign _6749 = _9338;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6751 <= _6748;
        else
            _6751 <= _6749;
    end
    assign _5661 = _6751;
    assign _5646 = _6625;
    assign _5647 = _6613;
    assign _5648 = _6597;
    assign _6587 = resetn & _6571;
    assign _6588 = _6587 & _5669;
    assign _5649 = _6588;
    assign _6589 = _5670 | _5666;
    assign _6590 = _6589 | _5668;
    assign _6571 = _6567 == _6570;
    assign _6591 = resetn & _6571;
    assign _6592 = _6591 & _6590;
    assign _5650 = _6592;
    assign _6618 = _5673[1:0];
    always @* begin
        case (_6618)
        0: _6619 <= _6614;
        1: _6619 <= _6615;
        2: _6619 <= _6616;
        default: _6619 <= _6617;
        endcase
    end
    assign _6622 = _5673[1:1];
    assign _6623 = _6622 ? _6621 : _6620;
    always @* begin
        case (_5667)
        0: _6625 <= _6624;
        1: _6625 <= _6623;
        default: _6625 <= _6619;
        endcase
    end
    assign _6701 = _6696 ? _6693 : _6625;
    assign _6702 = _6570 == _6567;
    assign _6703 = _6702 ? _6701 : _6688;
    assign _6686 = _6703;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6688 <= _6685;
        else
            _6688 <= _6686;
    end
    assign _5654 = _6688;
    assign _6609 = _5672[7:0];
    assign _6610 = { _6609, _6609 };
    assign _6611 = { _6610, _6610 };
    assign _6606 = _5672[15:0];
    assign _6607 = { _6606, _6606 };
    always @* begin
        case (_5667)
        0: _6613 <= _5672;
        1: _6613 <= _6607;
        default: _6613 <= _6611;
        endcase
    end
    assign _6704 = _6570 == _6567;
    assign _6705 = _6704 ? _6613 : _6684;
    assign _6682 = _6705;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6684 <= _6681;
        else
            _6684 <= _6682;
    end
    assign _5655 = _6684;
    assign _9390 = _7492 & _7484;
    assign _9391 = _9390 ? _7520 : _7507;
    assign _5674 = _9391;
    assign _6594 = _5673[31:2];
    assign _6595 = { _6594, _6593 };
    assign _6596 = _5666 | _5670;
    assign _6597 = _6596 ? _5674 : _6595;
    assign _6706 = _6570 == _6567;
    assign _6707 = _6706 ? _6597 : _6680;
    assign _6678 = _6707;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6680 <= _6677;
        else
            _6680 <= _6678;
    end
    assign _5656 = _6680;
    assign _6694 = _5666 | _5670;
    assign _6697 = _6696 ? _6694 : _6691;
    assign _6698 = _5669 ? gnd : _6697;
    assign _6699 = _6570 == _6567;
    assign _6700 = _6699 ? _6698 : _6691;
    assign _6689 = _6700;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6691 <= gnd;
        else
            _6691 <= _6689;
    end
    assign _5657 = _6691;
    assign _5658 = _6577;
    assign _9339 = _7683 ? _6743 : _6738;
    assign _9340 = _6763 ? _9339 : _6743;
    assign _9341 = _7696 ? _6743 : _9340;
    assign _9342 = _7789 ? _6743 : _9341;
    assign _9343 = _7920 ? _6740 : _6739;
    assign _9344 = _7464 ? _9343 : _6743;
    assign _9345 = _5634 ? _6740 : _9344;
    assign _9346 = vdd ? _9345 : _6737;
    assign _9347 = _7915 ? _6740 : _6739;
    assign _9348 = vdd ? _9346 : _9347;
    assign _9349 = _7826 ? _6735 : _6736;
    assign _9350 = _7828 ? _6734 : _9349;
    assign _9351 = vdd ? _9350 : _6737;
    assign _9352 = _7830 ? _6736 : _9351;
    assign _9353 = _7832 ? _6735 : _9352;
    assign _9354 = _7834 ? _6733 : _9353;
    assign _9355 = _7838 ? _6740 : _9354;
    assign _9356 = _7874 ? _6740 : _9355;
    assign _9357 = _7880 ? _6740 : _9356;
    assign _9358 = _7886 ? _6740 : _9357;
    assign _9359 = _7890 ? _6740 : _9358;
    assign _9360 = _7894 ? _6736 : _9359;
    assign _9361 = _7910 ? _6740 : _9360;
    assign _9362 = _7925 ? _9348 : _9361;
    assign _9363 = _7935 ? _6740 : _6739;
    assign _9364 = _7464 ? _9363 : _6743;
    assign _9365 = _5634 ? _6740 : _9364;
    assign _9366 = _7928 ? _6735 : _6736;
    assign _9367 = _7930 ? _6734 : _9366;
    assign _9368 = _7940 ? _9365 : _9367;
    assign _9369 = _5659 ? _6740 : _6743;
    assign _9370 = _7948 ? _9369 : _6740;
    assign _9371 = _8005 ? _6740 : _6743;
    assign _9372 = _8010 ? _6740 : _6743;
    assign _9373 = _8025 ? _9372 : _6743;
    assign _9374 = _8050 ? _6740 : _6743;
    assign _7674 = _5645[43:43];
    assign _7675 = ~ _7674;
    assign _7676 = _5645[3:3];
    assign _7677 = ~ _7676;
    assign _7678 = _7677 & _7675;
    assign _9288 = _7683 ? _6771 : _7678;
    assign _9289 = _6763 ? _9288 : _6771;
    assign _9290 = _7696 ? _6771 : _9289;
    assign _9291 = _7789 ? _6771 : _9290;
    assign _9292 = _6743 == _6740;
    assign _9293 = _9292 ? _9291 : _6771;
    assign _6572 = _6564 == _6570;
    assign _6581 = _6572 & _5670;
    assign _6582 = _5670 | _5668;
    assign _6583 = _6582 | _5669;
    assign _6718 = _6696 ? _6566 : _6570;
    assign _6719 = _5669 ? _6565 : _6718;
    assign _6692 = _5670 | _5668;
    assign _6720 = _6692 ? _6567 : _6564;
    assign _6721 = mem_ready ? _6720 : _6570;
    assign _6722 = mem_ready ? _6567 : _6570;
    assign _9174 = _7536[0:0];
    assign _9175 = _7536[1:1];
    assign _9176 = _7536[2:2];
    assign _9177 = _7536[3:3];
    assign _9178 = _7536[4:4];
    assign _9179 = _7536[5:5];
    assign _9180 = _7536[6:6];
    assign _9181 = _7536[7:7];
    assign _9182 = _7536[8:8];
    assign _9183 = _7536[9:9];
    assign _9184 = _7536[10:10];
    assign _9185 = _7536[11:11];
    assign _9186 = _7536[12:12];
    assign _9187 = _7536[13:13];
    assign _9188 = _7536[14:14];
    assign _9189 = _7536[15:15];
    assign _9190 = _7536[16:16];
    assign _9191 = _7536[17:17];
    assign _9192 = _7536[18:18];
    assign _9193 = _7536[19:19];
    assign _9194 = _7536[20:20];
    assign _9195 = _7536[21:21];
    assign _9196 = _7536[22:22];
    assign _9197 = _7536[23:23];
    assign _9198 = _7536[24:24];
    assign _9199 = _7536[25:25];
    assign _9200 = _7536[26:26];
    assign _9201 = _7536[27:27];
    assign _9202 = _7536[28:28];
    assign _9203 = _7536[29:29];
    assign _9204 = _7536[30:30];
    assign _9205 = _7536[31:31];
    assign _9206 = _9205 | _9204;
    assign _9207 = _9206 | _9203;
    assign _9208 = _9207 | _9202;
    assign _9209 = _9208 | _9201;
    assign _9210 = _9209 | _9200;
    assign _9211 = _9210 | _9199;
    assign _9212 = _9211 | _9198;
    assign _9213 = _9212 | _9197;
    assign _9214 = _9213 | _9196;
    assign _9215 = _9214 | _9195;
    assign _9216 = _9215 | _9194;
    assign _9217 = _9216 | _9193;
    assign _9218 = _9217 | _9192;
    assign _9219 = _9218 | _9191;
    assign _9220 = _9219 | _9190;
    assign _9221 = _9220 | _9189;
    assign _9222 = _9221 | _9188;
    assign _9223 = _9222 | _9187;
    assign _9224 = _9223 | _9186;
    assign _9225 = _9224 | _9185;
    assign _9226 = _9225 | _9184;
    assign _9227 = _9226 | _9183;
    assign _9228 = _9227 | _9182;
    assign _9229 = _9228 | _9181;
    assign _9230 = _9229 | _9180;
    assign _9231 = _9230 | _9179;
    assign _9232 = _9231 | _9178;
    assign _9233 = _9232 | _9177;
    assign _9234 = _9233 | _9176;
    assign _9235 = _9234 | _9175;
    assign _9236 = _9235 | _9174;
    assign _9237 = _9236 ? _7689 : _9173;
    assign _9238 = _7683 ? _7682 : _7679;
    assign _7813 = ~ _7472;
    assign _7814 = ~ _6763;
    assign _7815 = _7814 & _7813;
    assign _9171 = _7806 ? _7803 : _7815;
    assign _9172 = _7492 ? _7815 : _9171;
    assign _9173 = _7484 ? _7815 : _9172;
    assign _9239 = _6763 ? _9238 : _9173;
    assign _9240 = _7696 ? _9237 : _9239;
    assign _9241 = _7789 ? _9173 : _9240;
    assign _9242 = _5634 ? _7922 : _6787;
    assign _9243 = vdd ? _9242 : _6787;
    assign _9244 = vdd ? _9243 : _6787;
    assign _7826 = _5644[5:5];
    assign _9245 = _7826 ? _6787 : _6771;
    assign _7828 = _5644[4:4];
    assign _9246 = _7828 ? _7827 : _9245;
    assign _9247 = vdd ? _9246 : _6787;
    assign _9248 = _7830 ? _6771 : _9247;
    assign _9249 = _7832 ? _6787 : _9248;
    assign _9250 = _7834 ? _7833 : _9249;
    assign _9251 = _7838 ? _6787 : _9250;
    assign _9252 = _7874 ? _6787 : _9251;
    assign _9253 = _7880 ? _6787 : _9252;
    assign _9254 = _7886 ? _6787 : _9253;
    assign _9255 = _7890 ? _6787 : _9254;
    assign _9256 = _7894 ? _6771 : _9255;
    assign _9257 = _7910 ? _6787 : _9256;
    assign _9258 = _7925 ? _9244 : _9257;
    assign _9259 = _5634 ? _7937 : _6787;
    assign _7928 = _5644[5:5];
    assign _9260 = _7928 ? _6787 : _6771;
    assign _7930 = _5644[4:4];
    assign _9261 = _7930 ? _7929 : _9260;
    assign _9262 = _7940 ? _9259 : _9261;
    assign _9263 = _8005 ? _6771 : _6787;
    assign _9264 = _6743 == _6735;
    assign _9265 = _9264 ? _9263 : _6787;
    assign _9266 = _6743 == _6737;
    assign _9267 = _9266 ? _9262 : _9265;
    assign _9268 = _6743 == _6738;
    assign _9269 = _9268 ? _9258 : _9267;
    assign _9270 = _6743 == _6740;
    assign _9271 = _9270 ? _9241 : _9269;
    assign _9272 = _5659 ? _8079 : _9271;
    assign _8279 = _7422 ? _7945 : gnd;
    assign _6441 = _6308[2:2];
    assign _6440 = _6308[1:1];
    assign _6439 = _6308[0:0];
    assign _6442 = _6439 | _6440;
    assign _6443 = _6442 | _6441;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lui_auipc_jal <= gnd;
        else
            is_lui_auipc_jal <= _6443;
    end
    assign _6369 = _5652[31:25];
    assign _6371 = _6369 == _6370;
    assign _6372 = _5652[14:12];
    assign _6374 = _6372 == _6373;
    assign _6375 = _6374 & _6371;
    assign _6376 = _5652[31:25];
    assign _6378 = _6376 == _6377;
    assign _6379 = _5652[14:12];
    assign _6381 = _6379 == _6380;
    assign _6382 = _6381 & _6378;
    assign _6383 = _5652[31:25];
    assign _6385 = _6383 == _6384;
    assign _6386 = _5652[14:12];
    assign _6388 = _6386 == _6387;
    assign _6389 = _6388 & _6385;
    assign _6390 = _6389 | _6382;
    assign _6391 = _6390 | _6375;
    assign _6392 = is_alu_reg_imm & _6391;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_slli_srli_srai <= gnd;
        else
            if (_5846)
                is_slli_srli_srai <= _6392;
    end
    assign _6342 = _5652[14:12];
    assign _6344 = _6342 == _6343;
    assign _6345 = _5652[14:12];
    assign _6347 = _6345 == _6346;
    assign _6348 = _5652[14:12];
    assign _6350 = _6348 == _6349;
    assign _6351 = _5652[14:12];
    assign _6353 = _6351 == _6352;
    assign _6354 = _5652[14:12];
    assign _6356 = _6354 == _6355;
    assign _6357 = _5652[14:12];
    assign _6359 = _6357 == _6358;
    assign _6360 = _6359 | _6356;
    assign _6361 = _6360 | _6353;
    assign _6362 = _6361 | _6350;
    assign _6363 = _6362 | _6347;
    assign _6364 = _6363 | _6344;
    assign _6365 = is_alu_reg_imm & _6364;
    assign _6366 = instr_jalr | _6365;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_jalr_addi_slti_sltiu_xori_ori_andi <= gnd;
        else
            if (_5846)
                is_jalr_addi_slti_sltiu_xori_ori_andi <= _6366;
    end
    assign _6316 = _5652[31:25];
    assign _6318 = _6316 == _6317;
    assign _6319 = _5652[14:12];
    assign _6321 = _6319 == _6320;
    assign _6322 = _6321 & _6318;
    assign _6323 = _5652[31:25];
    assign _6325 = _6323 == _6324;
    assign _6326 = _5652[14:12];
    assign _6328 = _6326 == _6327;
    assign _6329 = _6328 & _6325;
    assign _6330 = _5652[31:25];
    assign _6332 = _6330 == _6331;
    assign _6333 = _5652[14:12];
    assign _6335 = _6333 == _6334;
    assign _6336 = _6335 & _6332;
    assign _6337 = _6336 | _6329;
    assign _6338 = _6337 | _6322;
    assign _6339 = is_alu_reg_reg & _6338;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sll_srl_sra <= gnd;
        else
            if (_5846)
                is_sll_srl_sra <= _6339;
    end
    assign _6431 = _6308[27:27];
    assign _6430 = _6308[18:18];
    assign _6429 = _6308[3:3];
    assign _6428 = _6308[2:2];
    assign _6427 = _6308[1:1];
    assign _6426 = _6308[0:0];
    assign _6432 = _6426 | _6427;
    assign _6433 = _6432 | _6428;
    assign _6434 = _6433 | _6429;
    assign _6435 = _6434 | _6430;
    assign _6436 = _6435 | _6431;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lui_auipc_jal_jalr_addi_add <= gnd;
        else
            is_lui_auipc_jal_jalr_addi_add <= _6436;
    end
    assign _6421 = _6308[30:30];
    assign _6420 = _6308[6:6];
    assign _6419 = _6308[19:19];
    assign _6422 = _6419 | _6420;
    assign _6423 = _6422 | _6421;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_slti_blt_slt <= gnd;
        else
            is_slti_blt_slt <= _6423;
    end
    assign _6414 = _6308[31:31];
    assign _6413 = _6308[8:8];
    assign _6412 = _6308[20:20];
    assign _6415 = _6412 | _6413;
    assign _6416 = _6415 | _6414;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sltiu_bltu_sltu <= gnd;
        else
            is_sltiu_bltu_sltu <= _6416;
    end
    assign _6407 = _6308[12:12];
    assign _6406 = _6308[14:14];
    assign _6405 = _6308[13:13];
    assign _6408 = _6405 | _6406;
    assign _6409 = _6408 | _6407;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lbu_lhu_lw <= gnd;
        else
            is_lbu_lhu_lw <= _6409;
    end
    assign _6398 = _6308[31:31];
    assign _6397 = _6308[20:20];
    assign _6396 = _6308[30:30];
    assign _6395 = _6308[19:19];
    assign _6399 = _6395 | _6396;
    assign _6400 = _6399 | _6397;
    assign _6401 = _6400 | _6398;
    assign _6402 = _6401 | is_beq_bne_blt_bge_bltu_bgeu;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_compare <= gnd;
        else
            is_compare <= _6402;
    end
    assign _6312 = _6308[40:40];
    assign _6311 = _6308[39:39];
    assign _6310 = _6308[38:38];
    assign _5892 = _5652[31:25];
    assign _5894 = _5892 == _5893;
    assign _5895 = _5652[6:0];
    assign _5897 = _5895 == _5896;
    assign _5898 = _5897 & _5894;
    assign _5899 = _5898 & vdd;
    assign _5900 = _5899 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_timer <= gnd;
        else
            if (_5846)
                instr_timer <= _5900;
    end
    assign _5903 = _5652[31:25];
    assign _5905 = _5903 == _5904;
    assign _5906 = _5652[6:0];
    assign _5908 = _5906 == _5907;
    assign _5909 = _5908 & _5905;
    assign _5910 = _5909 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_maskirq <= gnd;
        else
            if (_5846)
                instr_maskirq <= _5910;
    end
    assign _5913 = _5652[31:25];
    assign _5915 = _5913 == _5914;
    assign _5916 = _5652[6:0];
    assign _5918 = _5916 == _5917;
    assign _5919 = _5918 & _5915;
    assign _5920 = _5919 & vdd;
    assign _5921 = _5920 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_setq <= gnd;
        else
            if (_5846)
                instr_setq <= _5921;
    end
    assign _5924 = _5652[31:25];
    assign _5926 = _5924 == _5925;
    assign _5927 = _5652[6:0];
    assign _5929 = _5927 == _5928;
    assign _5930 = _5929 & _5926;
    assign _5931 = _5930 & vdd;
    assign _5932 = _5931 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_getq <= gnd;
        else
            if (_5846)
                instr_getq <= _5932;
    end
    assign _5935 = _5652[31:12];
    assign _5937 = _5935 == _5936;
    assign _5938 = _5652[6:0];
    assign _5940 = _5938 == _5939;
    assign _5941 = _5940 & _5937;
    assign _5942 = _5941 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdinstrh <= gnd;
        else
            if (_5846)
                instr_rdinstrh <= _5942;
    end
    assign _5945 = _5652[31:12];
    assign _5947 = _5945 == _5946;
    assign _5948 = _5652[6:0];
    assign _5950 = _5948 == _5949;
    assign _5951 = _5950 & _5947;
    assign _5952 = _5951 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdinstr <= gnd;
        else
            if (_5846)
                instr_rdinstr <= _5952;
    end
    assign _5955 = _5652[31:12];
    assign _5957 = _5955 == _5956;
    assign _5958 = _5652[6:0];
    assign _5960 = _5958 == _5959;
    assign _5961 = _5960 & _5957;
    assign _5962 = _5652[31:12];
    assign _5964 = _5962 == _5963;
    assign _5965 = _5652[6:0];
    assign _5967 = _5965 == _5966;
    assign _5968 = _5967 & _5964;
    assign _5969 = _5968 | _5961;
    assign _5970 = _5969 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdcycleh <= gnd;
        else
            if (_5846)
                instr_rdcycleh <= _5970;
    end
    assign _5973 = _5652[31:12];
    assign _5975 = _5973 == _5974;
    assign _5976 = _5652[6:0];
    assign _5978 = _5976 == _5977;
    assign _5979 = _5978 & _5975;
    assign _5980 = _5652[31:12];
    assign _5982 = _5980 == _5981;
    assign _5983 = _5652[6:0];
    assign _5985 = _5983 == _5984;
    assign _5986 = _5985 & _5982;
    assign _5987 = _5986 | _5979;
    assign _5988 = _5987 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdcycle <= gnd;
        else
            if (_5846)
                instr_rdcycle <= _5988;
    end
    assign _5991 = _5652[31:25];
    assign _5993 = _5991 == _5992;
    assign _5994 = _5652[14:12];
    assign _5996 = _5994 == _5995;
    assign _5997 = is_alu_reg_reg & _5996;
    assign _5998 = _5997 & _5993;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_and <= gnd;
        else
            if (_5846)
                instr_and <= _5998;
    end
    assign _6001 = _5652[31:25];
    assign _6003 = _6001 == _6002;
    assign _6004 = _5652[14:12];
    assign _6006 = _6004 == _6005;
    assign _6007 = is_alu_reg_reg & _6006;
    assign _6008 = _6007 & _6003;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_or <= gnd;
        else
            if (_5846)
                instr_or <= _6008;
    end
    assign _6011 = _5652[31:25];
    assign _6013 = _6011 == _6012;
    assign _6014 = _5652[14:12];
    assign _6016 = _6014 == _6015;
    assign _6017 = is_alu_reg_reg & _6016;
    assign _6018 = _6017 & _6013;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sra <= gnd;
        else
            if (_5846)
                instr_sra <= _6018;
    end
    assign _6021 = _5652[31:25];
    assign _6023 = _6021 == _6022;
    assign _6024 = _5652[14:12];
    assign _6026 = _6024 == _6025;
    assign _6027 = is_alu_reg_reg & _6026;
    assign _6028 = _6027 & _6023;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srl <= gnd;
        else
            if (_5846)
                instr_srl <= _6028;
    end
    assign _6031 = _5652[31:25];
    assign _6033 = _6031 == _6032;
    assign _6034 = _5652[14:12];
    assign _6036 = _6034 == _6035;
    assign _6037 = is_alu_reg_reg & _6036;
    assign _6038 = _6037 & _6033;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_xor <= gnd;
        else
            if (_5846)
                instr_xor <= _6038;
    end
    assign _6041 = _5652[31:25];
    assign _6043 = _6041 == _6042;
    assign _6044 = _5652[14:12];
    assign _6046 = _6044 == _6045;
    assign _6047 = is_alu_reg_reg & _6046;
    assign _6048 = _6047 & _6043;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sltu <= gnd;
        else
            if (_5846)
                instr_sltu <= _6048;
    end
    assign _6051 = _5652[31:25];
    assign _6053 = _6051 == _6052;
    assign _6054 = _5652[14:12];
    assign _6056 = _6054 == _6055;
    assign _6057 = is_alu_reg_reg & _6056;
    assign _6058 = _6057 & _6053;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slt <= gnd;
        else
            if (_5846)
                instr_slt <= _6058;
    end
    assign _6061 = _5652[31:25];
    assign _6063 = _6061 == _6062;
    assign _6064 = _5652[14:12];
    assign _6066 = _6064 == _6065;
    assign _6067 = is_alu_reg_reg & _6066;
    assign _6068 = _6067 & _6063;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sll <= gnd;
        else
            if (_5846)
                instr_sll <= _6068;
    end
    assign _6071 = _5652[31:25];
    assign _6073 = _6071 == _6072;
    assign _6074 = _5652[14:12];
    assign _6076 = _6074 == _6075;
    assign _6077 = is_alu_reg_reg & _6076;
    assign _6078 = _6077 & _6073;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sub <= gnd;
        else
            if (_5846)
                instr_sub <= _6078;
    end
    assign _6081 = _5652[31:25];
    assign _6083 = _6081 == _6082;
    assign _6084 = _5652[14:12];
    assign _6086 = _6084 == _6085;
    assign _5887 = _5653[6:0];
    assign _5889 = _5887 == _5888;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_alu_reg_reg <= gnd;
        else
            if (_5844)
                is_alu_reg_reg <= _5889;
    end
    assign _6087 = is_alu_reg_reg & _6086;
    assign _6088 = _6087 & _6083;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_add <= gnd;
        else
            if (_5846)
                instr_add <= _6088;
    end
    assign _6091 = _5652[31:25];
    assign _6093 = _6091 == _6092;
    assign _6094 = _5652[14:12];
    assign _6096 = _6094 == _6095;
    assign _6097 = is_alu_reg_imm & _6096;
    assign _6098 = _6097 & _6093;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srai <= gnd;
        else
            if (_5846)
                instr_srai <= _6098;
    end
    assign _6101 = _5652[31:25];
    assign _6103 = _6101 == _6102;
    assign _6104 = _5652[14:12];
    assign _6106 = _6104 == _6105;
    assign _6107 = is_alu_reg_imm & _6106;
    assign _6108 = _6107 & _6103;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srli <= gnd;
        else
            if (_5846)
                instr_srli <= _6108;
    end
    assign _6111 = _5652[31:25];
    assign _6113 = _6111 == _6112;
    assign _6114 = _5652[14:12];
    assign _6116 = _6114 == _6115;
    assign _6117 = is_alu_reg_imm & _6116;
    assign _6118 = _6117 & _6113;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slli <= gnd;
        else
            if (_5846)
                instr_slli <= _6118;
    end
    assign _6121 = _5652[14:12];
    assign _6123 = _6121 == _6122;
    assign _6124 = is_alu_reg_imm & _6123;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_andi <= gnd;
        else
            if (_5846)
                instr_andi <= _6124;
    end
    assign _6127 = _5652[14:12];
    assign _6129 = _6127 == _6128;
    assign _6130 = is_alu_reg_imm & _6129;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_ori <= gnd;
        else
            if (_5846)
                instr_ori <= _6130;
    end
    assign _6133 = _5652[14:12];
    assign _6135 = _6133 == _6134;
    assign _6136 = is_alu_reg_imm & _6135;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_xori <= gnd;
        else
            if (_5846)
                instr_xori <= _6136;
    end
    assign _6139 = _5652[14:12];
    assign _6141 = _6139 == _6140;
    assign _6142 = is_alu_reg_imm & _6141;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sltiu <= gnd;
        else
            if (_5846)
                instr_sltiu <= _6142;
    end
    assign _6145 = _5652[14:12];
    assign _6147 = _6145 == _6146;
    assign _6148 = is_alu_reg_imm & _6147;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slti <= gnd;
        else
            if (_5846)
                instr_slti <= _6148;
    end
    assign _6151 = _5652[14:12];
    assign _6153 = _6151 == _6152;
    assign _5882 = _5653[6:0];
    assign _5884 = _5882 == _5883;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_alu_reg_imm <= gnd;
        else
            if (_5844)
                is_alu_reg_imm <= _5884;
    end
    assign _6154 = is_alu_reg_imm & _6153;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_addi <= gnd;
        else
            if (_5846)
                instr_addi <= _6154;
    end
    assign _6157 = _5652[14:12];
    assign _6159 = _6157 == _6158;
    assign _6160 = is_sb_sh_sw & _6159;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sw <= gnd;
        else
            if (_5846)
                instr_sw <= _6160;
    end
    assign _6163 = _5652[14:12];
    assign _6165 = _6163 == _6164;
    assign _6166 = is_sb_sh_sw & _6165;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sh <= gnd;
        else
            if (_5846)
                instr_sh <= _6166;
    end
    assign _6169 = _5652[14:12];
    assign _6171 = _6169 == _6170;
    assign _5877 = _5653[6:0];
    assign _5879 = _5877 == _5878;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sb_sh_sw <= gnd;
        else
            if (_5844)
                is_sb_sh_sw <= _5879;
    end
    assign _6172 = is_sb_sh_sw & _6171;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sb <= gnd;
        else
            if (_5846)
                instr_sb <= _6172;
    end
    assign _6175 = _5652[14:12];
    assign _6177 = _6175 == _6176;
    assign _6178 = is_lb_lh_lw_lbu_lhu & _6177;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lhu <= gnd;
        else
            if (_5846)
                instr_lhu <= _6178;
    end
    assign _6181 = _5652[14:12];
    assign _6183 = _6181 == _6182;
    assign _6184 = is_lb_lh_lw_lbu_lhu & _6183;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lbu <= gnd;
        else
            if (_5846)
                instr_lbu <= _6184;
    end
    assign _6187 = _5652[14:12];
    assign _6189 = _6187 == _6188;
    assign _6190 = is_lb_lh_lw_lbu_lhu & _6189;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lw <= gnd;
        else
            if (_5846)
                instr_lw <= _6190;
    end
    assign _6193 = _5652[14:12];
    assign _6195 = _6193 == _6194;
    assign _6196 = is_lb_lh_lw_lbu_lhu & _6195;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lh <= gnd;
        else
            if (_5846)
                instr_lh <= _6196;
    end
    assign _6199 = _5652[14:12];
    assign _6201 = _6199 == _6200;
    assign _5872 = _5653[6:0];
    assign _5874 = _5872 == _5873;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lb_lh_lw_lbu_lhu <= gnd;
        else
            if (_5844)
                is_lb_lh_lw_lbu_lhu <= _5874;
    end
    assign _6202 = is_lb_lh_lw_lbu_lhu & _6201;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lb <= gnd;
        else
            if (_5846)
                instr_lb <= _6202;
    end
    assign _6205 = _5652[14:12];
    assign _6207 = _6205 == _6206;
    assign _6208 = is_beq_bne_blt_bge_bltu_bgeu & _6207;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bgeu <= gnd;
        else
            if (_5846)
                instr_bgeu <= _6208;
    end
    assign _6211 = _5652[14:12];
    assign _6213 = _6211 == _6212;
    assign _6214 = is_beq_bne_blt_bge_bltu_bgeu & _6213;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bltu <= gnd;
        else
            if (_5846)
                instr_bltu <= _6214;
    end
    assign _6217 = _5652[14:12];
    assign _6219 = _6217 == _6218;
    assign _6220 = is_beq_bne_blt_bge_bltu_bgeu & _6219;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bge <= gnd;
        else
            if (_5846)
                instr_bge <= _6220;
    end
    assign _6223 = _5652[14:12];
    assign _6225 = _6223 == _6224;
    assign _6226 = is_beq_bne_blt_bge_bltu_bgeu & _6225;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_blt <= gnd;
        else
            if (_5846)
                instr_blt <= _6226;
    end
    assign _6229 = _5652[14:12];
    assign _6231 = _6229 == _6230;
    assign _6232 = is_beq_bne_blt_bge_bltu_bgeu & _6231;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bne <= gnd;
        else
            if (_5846)
                instr_bne <= _6232;
    end
    assign _5845 = ~ _5662;
    assign _7412 = _6799 == _6795;
    assign _7409 = _6799 == _6795;
    assign _7410 = ~ _7409;
    assign _7418 = _7413 ? _7412 : _7410;
    assign _7398 = _6795[30:0];
    assign _7399 = _6795[31:31];
    assign _7400 = ~ _7399;
    assign _7401 = { _7400, _7398 };
    assign _7402 = _6799[30:0];
    assign _7403 = _6799[31:31];
    assign _7404 = ~ _7403;
    assign _7405 = { _7404, _7402 };
    assign _7406 = _7405 < _7401;
    assign _7407 = ~ _7406;
    assign _7395 = _6799 < _6795;
    assign _7396 = ~ _7395;
    assign _7416 = _7408 ? _7407 : _7396;
    assign _7420 = _7419 ? _7418 : _7416;
    assign _7385 = _6795[30:0];
    assign _7386 = _6795[31:31];
    assign _7387 = ~ _7386;
    assign _7388 = { _7387, _7385 };
    assign _7389 = _6799[30:0];
    assign _7390 = _6799[31:31];
    assign _7391 = ~ _7390;
    assign _7392 = { _7391, _7389 };
    assign _7393 = _7392 < _7388;
    assign _9128 = vdd ? _7820 : _7927;
    assign _7892 = _5645[0:0];
    assign _7893 = _7892 ? _7891 : _7510;
    assign _9129 = _7838 ? _7927 : _7820;
    assign _9130 = _7874 ? _7927 : _9129;
    assign _9131 = _7880 ? _7927 : _9130;
    assign _9132 = _7886 ? _7927 : _9131;
    assign _9133 = _7890 ? _7927 : _9132;
    assign _9134 = _7894 ? _7893 : _9133;
    assign _9135 = _7910 ? _7927 : _9134;
    assign _9136 = _7925 ? _9128 : _9135;
    assign _7992 = _6799[27:0];
    assign _7993 = { _7992, _7991 };
    assign _7985 = _6799[31:4];
    assign _7987 = { _7986, _7985 };
    assign _7997 = _7996 ? _7993 : _7987;
    assign _7976 = _6799[31:4];
    assign _7977 = _6799[31:31];
    assign _7978 = { _7977, _7977 };
    assign _7979 = { _7978, _7978 };
    assign _7981 = { _7979, _7976 };
    assign _7988 = _5645[33:33];
    assign _7989 = _5645[25:25];
    assign _7990 = _7989 | _7988;
    assign _7994 = _5645[29:29];
    assign _7995 = _5645[24:24];
    assign _7996 = _7995 | _7994;
    assign _7998 = _7996 | _7990;
    assign _7999 = _7998 ? _7997 : _7981;
    assign _7965 = _6799[30:0];
    assign _7966 = { _7965, _7964 };
    assign _7958 = _6799[31:1];
    assign _7960 = { _7959, _7958 };
    assign _7970 = _7969 ? _7966 : _7960;
    assign _7952 = _6799[31:1];
    assign _7953 = _6799[31:31];
    assign _7954 = { _7953, _7952 };
    assign _7961 = _5645[33:33];
    assign _7962 = _5645[25:25];
    assign _7963 = _7962 | _7961;
    assign _7967 = _5645[29:29];
    assign _7968 = _5645[24:24];
    assign _7969 = _7968 | _7967;
    assign _7971 = _7969 | _7963;
    assign _7972 = _7971 ? _7970 : _7954;
    assign _9137 = _8003 ? _7999 : _7972;
    assign _7923 = _7825[4:0];
    assign _8682 = vdd ? _7923 : _8266;
    assign _8683 = vdd ? _8682 : _8266;
    assign _7831 = _5640[4:0];
    assign _7829 = _7825[4:0];
    assign _8684 = vdd ? _7829 : _8266;
    assign _8685 = _7830 ? _8266 : _8684;
    assign _8686 = _7832 ? _7831 : _8685;
    assign _8687 = _7834 ? _8266 : _8686;
    assign _8688 = _7838 ? _8266 : _8687;
    assign _8689 = _7874 ? _8266 : _8688;
    assign _8690 = _7880 ? _8266 : _8689;
    assign _8691 = _7886 ? _8266 : _8690;
    assign _8692 = _7890 ? _8266 : _8691;
    assign _8693 = _7894 ? _8266 : _8692;
    assign _8694 = _7910 ? _8266 : _8693;
    assign _8695 = _7925 ? _8683 : _8694;
    assign _7201 = _7200[0:0];
    assign _7202 = _6810 & _7201;
    assign _7809 = _7510 + _7808;
    assign _9103 = vdd ? _7809 : _6808;
    assign _7807 = _7488 ? _7516 : _7520;
    assign _9104 = vdd ? _7807 : _6808;
    assign _7691 = _7512 + _7690;
    assign _8805 = _7536[0:0];
    assign _8806 = _7536[1:1];
    assign _8807 = _7536[2:2];
    assign _8808 = _7536[3:3];
    assign _8809 = _7536[4:4];
    assign _8810 = _7536[5:5];
    assign _8811 = _7536[6:6];
    assign _8812 = _7536[7:7];
    assign _8813 = _7536[8:8];
    assign _8814 = _7536[9:9];
    assign _8815 = _7536[10:10];
    assign _8816 = _7536[11:11];
    assign _8817 = _7536[12:12];
    assign _8818 = _7536[13:13];
    assign _8819 = _7536[14:14];
    assign _8820 = _7536[15:15];
    assign _8821 = _7536[16:16];
    assign _8822 = _7536[17:17];
    assign _8823 = _7536[18:18];
    assign _8824 = _7536[19:19];
    assign _8825 = _7536[20:20];
    assign _8826 = _7536[21:21];
    assign _8827 = _7536[22:22];
    assign _8828 = _7536[23:23];
    assign _8829 = _7536[24:24];
    assign _8830 = _7536[25:25];
    assign _8831 = _7536[26:26];
    assign _8832 = _7536[27:27];
    assign _8833 = _7536[28:28];
    assign _8834 = _7536[29:29];
    assign _8835 = _7536[30:30];
    assign _8836 = _7536[31:31];
    assign _8837 = _8836 | _8835;
    assign _8838 = _8837 | _8834;
    assign _8839 = _8838 | _8833;
    assign _8840 = _8839 | _8832;
    assign _8841 = _8840 | _8831;
    assign _8842 = _8841 | _8830;
    assign _8843 = _8842 | _8829;
    assign _8844 = _8843 | _8828;
    assign _8845 = _8844 | _8827;
    assign _8846 = _8845 | _8826;
    assign _8847 = _8846 | _8825;
    assign _8848 = _8847 | _8824;
    assign _8849 = _8848 | _8823;
    assign _8850 = _8849 | _8822;
    assign _8851 = _8850 | _8821;
    assign _8852 = _8851 | _8820;
    assign _8853 = _8852 | _8819;
    assign _8854 = _8853 | _8818;
    assign _8855 = _8854 | _8817;
    assign _8856 = _8855 | _8816;
    assign _8857 = _8856 | _8815;
    assign _8858 = _8857 | _8814;
    assign _8859 = _8858 | _8813;
    assign _8860 = _8859 | _8812;
    assign _8861 = _8860 | _8811;
    assign _8862 = _8861 | _8810;
    assign _8863 = _8862 | _8809;
    assign _8864 = _8863 | _8808;
    assign _8865 = _8864 | _8807;
    assign _8866 = _8865 | _8806;
    assign _8867 = _8866 | _8805;
    assign _8868 = _8867 ? _7691 : _7512;
    assign _5638 = _6489;
    assign _7681 = _7512 + _5638;
    assign _7687 = _7512 + _7686;
    assign _8869 = _7683 ? _7681 : _7687;
    assign _7449 = _6799 + _6795;
    assign _7447 = _6799 - _6795;
    assign _7455 = _7450 ? _7449 : _7447;
    assign _7445 = { _7443, _7422 };
    assign _7432 = _6799 ^ _6795;
    assign _7453 = _7446 ? _7445 : _7432;
    assign _7457 = _7456 ? _7455 : _7453;
    assign _7428 = _6799 | _6795;
    assign _7424 = _6799 & _6795;
    assign _7429 = _5645[35:35];
    assign _7430 = _5645[22:22];
    assign _7431 = _7430 | _7429;
    assign _7451 = _7431 ? _7428 : _7424;
    assign _7433 = _5645[32:32];
    assign _7434 = _5645[21:21];
    assign _7435 = _7434 | _7433;
    assign _7446 = _5644[13:13];
    assign _7454 = _7446 | _7435;
    assign _7448 = _5645[28:28];
    assign _7450 = _5644[6:6];
    assign _7456 = _7450 | _7448;
    assign _7458 = _7456 | _7454;
    assign _7459 = _7458 ? _7457 : _7451;
    assign _7514 = _7459;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7516 <= _7513;
        else
            _7516 <= _7514;
    end
    assign _8704 = _7536[0:0];
    assign _8705 = _7536[1:1];
    assign _8706 = _7536[2:2];
    assign _8707 = _7536[3:3];
    assign _8708 = _7536[4:4];
    assign _8709 = _7536[5:5];
    assign _8710 = _7536[6:6];
    assign _8711 = _7536[7:7];
    assign _8712 = _7536[8:8];
    assign _8713 = _7536[9:9];
    assign _8714 = _7536[10:10];
    assign _8715 = _7536[11:11];
    assign _8716 = _7536[12:12];
    assign _8717 = _7536[13:13];
    assign _8718 = _7536[14:14];
    assign _8719 = _7536[15:15];
    assign _8720 = _7536[16:16];
    assign _8721 = _7536[17:17];
    assign _8722 = _7536[18:18];
    assign _8723 = _7536[19:19];
    assign _8724 = _7536[20:20];
    assign _8725 = _7536[21:21];
    assign _8726 = _7536[22:22];
    assign _8727 = _7536[23:23];
    assign _8728 = _7536[24:24];
    assign _8729 = _7536[25:25];
    assign _8730 = _7536[26:26];
    assign _8731 = _7536[27:27];
    assign _8732 = _7536[28:28];
    assign _8733 = _7536[29:29];
    assign _8734 = _7536[30:30];
    assign _8735 = _7536[31:31];
    assign _8736 = _8735 | _8734;
    assign _8737 = _8736 | _8733;
    assign _8738 = _8737 | _8732;
    assign _8739 = _8738 | _8731;
    assign _8740 = _8739 | _8730;
    assign _8741 = _8740 | _8729;
    assign _8742 = _8741 | _8728;
    assign _8743 = _8742 | _8727;
    assign _8744 = _8743 | _8726;
    assign _8745 = _8744 | _8725;
    assign _8746 = _8745 | _8724;
    assign _8747 = _8746 | _8723;
    assign _8748 = _8747 | _8722;
    assign _8749 = _8748 | _8721;
    assign _8750 = _8749 | _8720;
    assign _8751 = _8750 | _8719;
    assign _8752 = _8751 | _8718;
    assign _8753 = _8752 | _8717;
    assign _8754 = _8753 | _8716;
    assign _8755 = _8754 | _8715;
    assign _8756 = _8755 | _8714;
    assign _8757 = _8756 | _8713;
    assign _8758 = _8757 | _8712;
    assign _8759 = _8758 | _8711;
    assign _8760 = _8759 | _8710;
    assign _8761 = _8760 | _8709;
    assign _8762 = _8761 | _8708;
    assign _8763 = _8762 | _8707;
    assign _8764 = _8763 | _8706;
    assign _8765 = _8764 | _8705;
    assign _8766 = _8765 | _8704;
    assign _8767 = _8766 ? _7536 : _8265;
    assign _8768 = _7696 ? _8767 : _8265;
    assign _8769 = _7789 ? _8265 : _8768;
    assign _8770 = _5634 ? _5636 : _8265;
    assign _8771 = vdd ? _8770 : _8265;
    assign _8772 = vdd ? _8771 : _8265;
    assign _7902 = count_cycle[31:0];
    assign _8097 = count_cycle + _8096;
    assign _9007 = vdd ? _8097 : count_cycle;
    assign _7478 = _9007;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            count_cycle <= _7477;
        else
            count_cycle <= _7478;
    end
    assign _7900 = count_cycle[63:32];
    assign _7906 = _7903 ? _7902 : _7900;
    assign _7898 = _7476[31:0];
    assign _7685 = _7476 + _7684;
    assign _9008 = vdd ? _7685 : _7476;
    assign _9009 = _6763 ? _9008 : _7476;
    assign _9010 = _7696 ? _7476 : _9009;
    assign _9011 = _7789 ? _7476 : _9010;
    assign _9012 = _6743 == _6740;
    assign _9013 = _9012 ? _9011 : _7476;
    assign _7474 = _9013;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7476 <= _7473;
        else
            _7476 <= _7474;
    end
    assign _7896 = _7476[63:32];
    assign _7899 = _5645[39:39];
    assign _7904 = _7899 ? _7898 : _7896;
    assign _7901 = _5645[38:38];
    assign _7903 = _5645[37:37];
    assign _7907 = _7903 | _7901;
    assign _7908 = _7907 ? _7906 : _7904;
    assign _8773 = _7838 ? _7673 : _8265;
    assign _8774 = _7874 ? _7666 : _8773;
    assign _8775 = _7880 ? _7382 : _8774;
    assign _8776 = _7886 ? _7382 : _8775;
    assign _8777 = _7890 ? _7382 : _8776;
    assign _8778 = _7894 ? _8265 : _8777;
    assign _8779 = _7910 ? _7908 : _8778;
    assign _8780 = _7925 ? _8772 : _8779;
    assign _5825 = _5739[63:32];
    assign _5741 = _5740 ^ _5727;
    assign _5745 = _5735 & _5727;
    assign _5786 = _5672[31:31];
    assign _5787 = { _5786, _5786 };
    assign _5788 = { _5787, _5787 };
    assign _5789 = { _5788, _5788 };
    assign _5790 = { _5789, _5789 };
    assign _5791 = { _5790, _5790 };
    assign _5793 = { _5791, _5672 };
    assign _9151 = vdd ? _7825 : _7926;
    assign _9152 = vdd ? _9151 : _7926;
    assign _9153 = vdd ? _7825 : _7926;
    assign _7830 = _5644[3:3];
    assign _9154 = _7830 ? _5639 : _9153;
    assign _7832 = _5644[2:2];
    assign _9155 = _7832 ? _7926 : _9154;
    assign _7834 = _5644[1:1];
    assign _9156 = _7834 ? _7926 : _9155;
    assign _9157 = _7838 ? _7926 : _9156;
    assign _9158 = _7874 ? _7926 : _9157;
    assign _9159 = _7880 ? _7926 : _9158;
    assign _9160 = _7886 ? _7926 : _9159;
    assign _9161 = _7890 ? _7926 : _9160;
    assign _9162 = _7894 ? _5639 : _9161;
    assign _9163 = _7910 ? _7926 : _9162;
    assign _9164 = _7925 ? _9152 : _9163;
    assign _9165 = _6743 == _6737;
    assign _9166 = _9165 ? _7825 : _6795;
    assign _9167 = _6743 == _6738;
    assign _9168 = _9167 ? _9164 : _9166;
    assign _6793 = _9168;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6795 <= _6792;
        else
            _6795 <= _6793;
    end
    assign _5672 = _6795;
    assign _5785 = { _5783, _5672 };
    assign _5794 = _5699 ? _5793 : _5785;
    assign _5758 = _5727[62:0];
    assign _5759 = { _5758, _5757 };
    assign _5819 = _5766 ? _5794 : _5759;
    assign _5725 = _5819;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5727 <= _5724;
        else
            _5727 <= _5725;
    end
    assign _5746 = _5739 & _5727;
    assign _5747 = _5744 | _5746;
    assign _5748 = _5747 | _5745;
    assign _5744 = _5739 & _5735;
    assign _5749 = _5731[0:0];
    assign _5750 = _5749 ? _5748 : _5744;
    assign _5752 = _5750[62:0];
    assign _5753 = { _5752, _5751 };
    assign _5817 = _5766 ? _5777 : _5753;
    assign _5733 = _5817;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5735 <= _5732;
        else
            _5735 <= _5733;
    end
    assign _5740 = _5739 ^ _5735;
    assign _5802 = _5673[31:31];
    assign _5803 = { _5802, _5802 };
    assign _5804 = { _5803, _5803 };
    assign _5805 = { _5804, _5804 };
    assign _5806 = { _5805, _5805 };
    assign _5807 = { _5806, _5806 };
    assign _5809 = { _5807, _5673 };
    assign _5801 = { _5799, _5673 };
    assign _5717 = _5699 | _5705;
    assign _5810 = _5717 ? _5809 : _5801;
    assign _5754 = _5731[63:1];
    assign _5756 = { _5755, _5754 };
    assign _5818 = _5766 ? _5810 : _5756;
    assign _5729 = _5818;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5731 <= _5728;
        else
            _5731 <= _5729;
    end
    assign _5742 = _5731[0:0];
    assign _5743 = _5742 ? _5741 : _5740;
    assign _5816 = _5766 ? _5778 : _5743;
    assign _5737 = _5816;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5739 <= _5736;
        else
            _5739 <= _5737;
    end
    assign _5824 = _5739[31:0];
    assign _5826 = _5716 ? _5825 : _5824;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5829 <= _5827;
        else
            if (_5769)
                _5829 <= _5826;
    end
    assign _5839 = _5833 ? _5829 : _5838;
    assign _5840 = _5834 ? pcpi_rd : _5839;
    assign _5636 = _5840;
    assign _8781 = _5634 ? _5636 : _8265;
    assign _8782 = _7940 ? _8781 : _8265;
    assign _8803 = _6743 == _6740;
    assign _8804 = _8803 ? _7512 : _7510;
    assign _7508 = _8804;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7510 <= _39;
        else
            _7510 <= _7508;
    end
    assign _7949 = _7510 + _5639;
    assign _8783 = _8005 ? _6799 : _8265;
    assign _8037 = _5651[15:0];
    assign _8038 = _8037[15:15];
    assign _8039 = { _8038, _8038 };
    assign _8040 = { _8039, _8039 };
    assign _8041 = { _8040, _8040 };
    assign _8042 = { _8041, _8041 };
    assign _8044 = { _8042, _8037 };
    assign _8045 = _7504 ? _5651 : _8044;
    assign _6650 = mem_rdata[31:24];
    assign _6657 = { _6655, _6650 };
    assign _6642 = mem_rdata[23:16];
    assign _6649 = { _6647, _6642 };
    assign _6634 = mem_rdata[15:8];
    assign _6641 = { _6639, _6634 };
    assign _6626 = mem_rdata[7:0];
    assign _6633 = { _6631, _6626 };
    assign _6658 = _5673[1:0];
    always @* begin
        case (_6658)
        0: _6659 <= _6633;
        1: _6659 <= _6641;
        2: _6659 <= _6649;
        default: _6659 <= _6657;
        endcase
    end
    assign _6660 = mem_rdata[31:16];
    assign _6666 = { _6664, _6660 };
    assign _6667 = mem_rdata[15:0];
    assign _6673 = { _6671, _6667 };
    assign _5673 = _6799;
    assign _6674 = _5673[1:1];
    assign _6675 = _6674 ? _6666 : _6673;
    assign _8019 = _8018 ? _8017 : _8015;
    assign _8016 = _5645[16:16];
    assign _8018 = _5645[15:15];
    assign _8020 = _8018 | _8016;
    assign _8021 = _8020 ? _8019 : _8013;
    assign _9278 = _8023 ? _8021 : _6775;
    assign _9279 = _8025 ? _9278 : _6775;
    assign _8066 = _8065 ? _8062 : _8058;
    assign _8059 = _5645[14:14];
    assign _8060 = _5645[11:11];
    assign _8061 = _8060 | _8059;
    assign _8063 = _5645[13:13];
    assign _8064 = _5645[10:10];
    assign _8065 = _8064 | _8063;
    assign _8067 = _8065 | _8061;
    assign _8068 = _8067 ? _8066 : _8056;
    assign _9280 = _8070 ? _8068 : _6775;
    assign _9281 = _8072 ? _9280 : _6775;
    assign _9282 = _6743 == _6733;
    assign _9283 = _9282 ? _9281 : _6775;
    assign _9284 = _6743 == _6734;
    assign _9285 = _9284 ? _9279 : _9283;
    assign _9286 = _6743 == _6740;
    assign _9287 = _9286 ? _7812 : _9285;
    assign _6773 = _9287;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6775 <= _6772;
        else
            _6775 <= _6773;
    end
    assign _5667 = _6775;
    always @* begin
        case (_5667)
        0: _6676 <= mem_rdata;
        1: _6676 <= _6675;
        default: _6676 <= _6659;
        endcase
    end
    assign _5651 = _6676;
    assign _8028 = _5651[7:0];
    assign _8029 = _8028[7:7];
    assign _8030 = { _8029, _8029 };
    assign _8031 = { _8030, _8030 };
    assign _8032 = { _8031, _8031 };
    assign _8033 = { _8032, _8032 };
    assign _8034 = { _8033, _8032 };
    assign _8036 = { _8034, _8028 };
    assign _8054 = _5645[11:11];
    assign _8881 = _8070 ? _8054 : _7500;
    assign _8882 = _8072 ? _8881 : _7500;
    assign _8883 = _6743 == _6733;
    assign _8884 = _8883 ? _8882 : _7500;
    assign _8885 = _6743 == _6740;
    assign _8886 = _8885 ? _7791 : _8884;
    assign _7498 = _8886;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7500 <= _7497;
        else
            _7500 <= _7498;
    end
    assign _8055 = _5644[10:10];
    assign _8875 = _8070 ? _8055 : _7504;
    assign _8876 = _8072 ? _8875 : _7504;
    assign _8877 = _6743 == _6733;
    assign _8878 = _8877 ? _8876 : _7504;
    assign _8879 = _6743 == _6740;
    assign _8880 = _8879 ? _7792 : _8878;
    assign _7502 = _8880;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7504 <= _7501;
        else
            _7504 <= _7502;
    end
    assign _8046 = _7504 | _7500;
    assign _8047 = _8046 ? _8045 : _8036;
    assign _8784 = _8050 ? _8047 : _8265;
    assign _8785 = _8072 ? _8784 : _8265;
    assign _8786 = _6743 == _6733;
    assign _8787 = _8786 ? _8785 : _8265;
    assign _8788 = _6743 == _6735;
    assign _8789 = _8788 ? _8783 : _8787;
    assign _8790 = _6743 == _6736;
    assign _8791 = _8790 ? _7949 : _8789;
    assign _8792 = _6743 == _6737;
    assign _8793 = _8792 ? _8782 : _8791;
    assign _8794 = _6743 == _6738;
    assign _8795 = _8794 ? _8780 : _8793;
    assign _8796 = _6743 == _6740;
    assign _8797 = _8796 ? _8769 : _8795;
    assign _7518 = _8797;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7520 <= _7517;
        else
            _7520 <= _7518;
    end
    assign _8985 = _7948 ? _7488 : _7942;
    assign _8986 = _6743 == _6736;
    assign _8987 = _8986 ? _8985 : _7488;
    assign _8988 = _6743 == _6740;
    assign _8989 = _8988 ? _7794 : _8987;
    assign _7486 = _8989;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7488 <= _7485;
        else
            _7488 <= _7486;
    end
    assign _7810 = _7488 ? _7516 : _7520;
    assign _7811 = _7492 ? _7810 : _7507;
    assign _8798 = _7806 ? _40 : _7507;
    assign _8799 = _7492 ? _7507 : _8798;
    assign _8800 = _7484 ? _7811 : _8799;
    assign _8801 = _6743 == _6740;
    assign _8802 = _8801 ? _8800 : _7511;
    assign _7512 = _8802;
    assign _8870 = _6763 ? _8869 : _7512;
    assign _8871 = _7696 ? _8868 : _8870;
    assign _8872 = _7789 ? _7512 : _8871;
    assign _8873 = _6743 == _6740;
    assign _8874 = _8873 ? _8872 : _7507;
    assign _7505 = _8874;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7507 <= _39;
        else
            _7507 <= _7505;
    end
    assign _9105 = vdd ? _7507 : _6808;
    assign _7797 = ~ _7666;
    assign _7798 = _7536 & _7797;
    assign _9106 = vdd ? _7798 : _6808;
    assign _9107 = _7802 ? _9106 : _6808;
    assign _9108 = _7806 ? _9105 : _9107;
    assign _9109 = _7492 ? _9104 : _9108;
    assign _7683 = _5645[2:2];
    assign _8990 = _7683 ? _7680 : _7793;
    assign _8991 = _6763 ? _8990 : _7793;
    assign _8992 = _7696 ? _7793 : _8991;
    assign _7717 = _7528[0:0];
    assign _7718 = _7528[1:1];
    assign _7719 = _7718 | _7717;
    assign _7722 = _7721[0:0];
    assign _7723 = _7721[1:1];
    assign _7724 = _7721[2:2];
    assign _7725 = _7721[3:3];
    assign _7726 = _7721[4:4];
    assign _7727 = _7721[5:5];
    assign _7728 = _7721[6:6];
    assign _7729 = _7721[7:7];
    assign _7730 = _7721[8:8];
    assign _7731 = _7721[9:9];
    assign _7732 = _7721[10:10];
    assign _7733 = _7721[11:11];
    assign _7734 = _7721[12:12];
    assign _7735 = _7721[13:13];
    assign _7736 = _7721[14:14];
    assign _7737 = _7721[15:15];
    assign _7738 = _7721[16:16];
    assign _7739 = _7721[17:17];
    assign _7740 = _7721[18:18];
    assign _7741 = _7721[19:19];
    assign _7742 = _7721[20:20];
    assign _7743 = _7721[21:21];
    assign _7744 = _7721[22:22];
    assign _7745 = _7721[23:23];
    assign _7746 = _7721[24:24];
    assign _7747 = _7721[25:25];
    assign _7748 = _7721[26:26];
    assign _7749 = _7721[27:27];
    assign _7750 = _7721[28:28];
    assign _7751 = _7721[29:29];
    assign _7752 = _7721[30:30];
    assign _7720 = ~ _7666;
    assign _7721 = _7536 & _7720;
    assign _7753 = _7721[31:31];
    assign _7754 = _7753 | _7752;
    assign _7755 = _7754 | _7751;
    assign _7756 = _7755 | _7750;
    assign _7757 = _7756 | _7749;
    assign _7758 = _7757 | _7748;
    assign _7759 = _7758 | _7747;
    assign _7760 = _7759 | _7746;
    assign _7761 = _7760 | _7745;
    assign _7762 = _7761 | _7744;
    assign _7763 = _7762 | _7743;
    assign _7764 = _7763 | _7742;
    assign _7765 = _7764 | _7741;
    assign _7766 = _7765 | _7740;
    assign _7767 = _7766 | _7739;
    assign _7768 = _7767 | _7738;
    assign _7769 = _7768 | _7737;
    assign _7770 = _7769 | _7736;
    assign _7771 = _7770 | _7735;
    assign _7772 = _7771 | _7734;
    assign _7773 = _7772 | _7733;
    assign _7774 = _7773 | _7732;
    assign _7775 = _7774 | _7731;
    assign _7776 = _7775 | _7730;
    assign _7777 = _7776 | _7729;
    assign _7778 = _7777 | _7728;
    assign _7779 = _7778 | _7727;
    assign _7780 = _7779 | _7726;
    assign _7781 = _7780 | _7725;
    assign _7782 = _7781 | _7724;
    assign _7783 = _7782 | _7723;
    assign _7784 = _7783 | _7722;
    assign _8666 = _7806 ? _7804 : _7532;
    assign _8893 = _7536[0:0];
    assign _8894 = _7536[1:1];
    assign _8895 = _7536[2:2];
    assign _8896 = _7536[3:3];
    assign _8897 = _7536[4:4];
    assign _8898 = _7536[5:5];
    assign _8899 = _7536[6:6];
    assign _8900 = _7536[7:7];
    assign _8901 = _7536[8:8];
    assign _8902 = _7536[9:9];
    assign _8903 = _7536[10:10];
    assign _8904 = _7536[11:11];
    assign _8905 = _7536[12:12];
    assign _8906 = _7536[13:13];
    assign _8907 = _7536[14:14];
    assign _8908 = _7536[15:15];
    assign _8909 = _7536[16:16];
    assign _8910 = _7536[17:17];
    assign _8911 = _7536[18:18];
    assign _8912 = _7536[19:19];
    assign _8913 = _7536[20:20];
    assign _8914 = _7536[21:21];
    assign _8915 = _7536[22:22];
    assign _8916 = _7536[23:23];
    assign _8917 = _7536[24:24];
    assign _8918 = _7536[25:25];
    assign _8919 = _7536[26:26];
    assign _8920 = _7536[27:27];
    assign _8921 = _7536[28:28];
    assign _8922 = _7536[29:29];
    assign _8923 = _7536[30:30];
    assign _8924 = _7536[31:31];
    assign _8925 = _8924 | _8923;
    assign _8926 = _8925 | _8922;
    assign _8927 = _8926 | _8921;
    assign _8928 = _8927 | _8920;
    assign _8929 = _8928 | _8919;
    assign _8930 = _8929 | _8918;
    assign _8931 = _8930 | _8917;
    assign _8932 = _8931 | _8916;
    assign _8933 = _8932 | _8915;
    assign _8934 = _8933 | _8914;
    assign _8935 = _8934 | _8913;
    assign _8936 = _8935 | _8912;
    assign _8937 = _8936 | _8911;
    assign _8938 = _8937 | _8910;
    assign _8939 = _8938 | _8909;
    assign _8940 = _8939 | _8908;
    assign _8941 = _8940 | _8907;
    assign _8942 = _8941 | _8906;
    assign _8943 = _8942 | _8905;
    assign _8944 = _8943 | _8904;
    assign _8945 = _8944 | _8903;
    assign _8946 = _8945 | _8902;
    assign _8947 = _8946 | _8901;
    assign _8948 = _8947 | _8900;
    assign _8949 = _8948 | _8899;
    assign _8950 = _8949 | _8898;
    assign _8951 = _8950 | _8897;
    assign _8952 = _8951 | _8896;
    assign _8953 = _8952 | _8895;
    assign _8954 = _8953 | _8894;
    assign _8955 = _8954 | _8893;
    assign _8956 = _8955 ? _7692 : _7795;
    assign _7693 = _5645[45:45];
    assign _9014 = _7536[0:0];
    assign _9015 = _7536[1:1];
    assign _9016 = _7536[2:2];
    assign _9017 = _7536[3:3];
    assign _9018 = _7536[4:4];
    assign _9019 = _7536[5:5];
    assign _9020 = _7536[6:6];
    assign _9021 = _7536[7:7];
    assign _9022 = _7536[8:8];
    assign _9023 = _7536[9:9];
    assign _9024 = _7536[10:10];
    assign _9025 = _7536[11:11];
    assign _9026 = _7536[12:12];
    assign _9027 = _7536[13:13];
    assign _9028 = _7536[14:14];
    assign _9029 = _7536[15:15];
    assign _9030 = _7536[16:16];
    assign _9031 = _7536[17:17];
    assign _9032 = _7536[18:18];
    assign _9033 = _7536[19:19];
    assign _9034 = _7536[20:20];
    assign _9035 = _7536[21:21];
    assign _9036 = _7536[22:22];
    assign _9037 = _7536[23:23];
    assign _9038 = _7536[24:24];
    assign _9039 = _7536[25:25];
    assign _9040 = _7536[26:26];
    assign _9041 = _7536[27:27];
    assign _9042 = _7536[28:28];
    assign _9043 = _7536[29:29];
    assign _9044 = _7536[30:30];
    assign _7840 = _7839[0:0];
    assign _8601 = vdd ? _7840 : _7572;
    assign _8602 = _7874 ? _8601 : _7572;
    assign _8603 = _7880 ? _7572 : _8602;
    assign _8604 = _7886 ? _7572 : _8603;
    assign _8605 = _7890 ? _7572 : _8604;
    assign _8606 = _7894 ? _7572 : _8605;
    assign _8607 = _7910 ? _7572 : _8606;
    assign _8608 = _7925 ? _7572 : _8607;
    assign _8609 = _6743 == _6738;
    assign _8610 = _8609 ? _8608 : _7572;
    assign _7570 = _8610;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7572 <= vdd;
        else
            _7572 <= _7570;
    end
    assign _7842 = _7839[2:2];
    assign _8581 = vdd ? _7842 : _7578;
    assign _8582 = _7874 ? _8581 : _7578;
    assign _8583 = _7880 ? _7578 : _8582;
    assign _8584 = _7886 ? _7578 : _8583;
    assign _8585 = _7890 ? _7578 : _8584;
    assign _8586 = _7894 ? _7578 : _8585;
    assign _8587 = _7910 ? _7578 : _8586;
    assign _8588 = _7925 ? _7578 : _8587;
    assign _8589 = _6743 == _6738;
    assign _8590 = _8589 ? _8588 : _7578;
    assign _7576 = _8590;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7578 <= vdd;
        else
            _7578 <= _7576;
    end
    assign _7843 = _7839[3:3];
    assign _8571 = vdd ? _7843 : _7581;
    assign _8572 = _7874 ? _8571 : _7581;
    assign _8573 = _7880 ? _7581 : _8572;
    assign _8574 = _7886 ? _7581 : _8573;
    assign _8575 = _7890 ? _7581 : _8574;
    assign _8576 = _7894 ? _7581 : _8575;
    assign _8577 = _7910 ? _7581 : _8576;
    assign _8578 = _7925 ? _7581 : _8577;
    assign _8579 = _6743 == _6738;
    assign _8580 = _8579 ? _8578 : _7581;
    assign _7579 = _8580;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7581 <= vdd;
        else
            _7581 <= _7579;
    end
    assign _7844 = _7839[4:4];
    assign _8561 = vdd ? _7844 : _7584;
    assign _8562 = _7874 ? _8561 : _7584;
    assign _8563 = _7880 ? _7584 : _8562;
    assign _8564 = _7886 ? _7584 : _8563;
    assign _8565 = _7890 ? _7584 : _8564;
    assign _8566 = _7894 ? _7584 : _8565;
    assign _8567 = _7910 ? _7584 : _8566;
    assign _8568 = _7925 ? _7584 : _8567;
    assign _8569 = _6743 == _6738;
    assign _8570 = _8569 ? _8568 : _7584;
    assign _7582 = _8570;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7584 <= vdd;
        else
            _7584 <= _7582;
    end
    assign _7845 = _7839[5:5];
    assign _8551 = vdd ? _7845 : _7587;
    assign _8552 = _7874 ? _8551 : _7587;
    assign _8553 = _7880 ? _7587 : _8552;
    assign _8554 = _7886 ? _7587 : _8553;
    assign _8555 = _7890 ? _7587 : _8554;
    assign _8556 = _7894 ? _7587 : _8555;
    assign _8557 = _7910 ? _7587 : _8556;
    assign _8558 = _7925 ? _7587 : _8557;
    assign _8559 = _6743 == _6738;
    assign _8560 = _8559 ? _8558 : _7587;
    assign _7585 = _8560;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7587 <= vdd;
        else
            _7587 <= _7585;
    end
    assign _7846 = _7839[6:6];
    assign _8541 = vdd ? _7846 : _7590;
    assign _8542 = _7874 ? _8541 : _7590;
    assign _8543 = _7880 ? _7590 : _8542;
    assign _8544 = _7886 ? _7590 : _8543;
    assign _8545 = _7890 ? _7590 : _8544;
    assign _8546 = _7894 ? _7590 : _8545;
    assign _8547 = _7910 ? _7590 : _8546;
    assign _8548 = _7925 ? _7590 : _8547;
    assign _8549 = _6743 == _6738;
    assign _8550 = _8549 ? _8548 : _7590;
    assign _7588 = _8550;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7590 <= vdd;
        else
            _7590 <= _7588;
    end
    assign _7847 = _7839[7:7];
    assign _8531 = vdd ? _7847 : _7593;
    assign _8532 = _7874 ? _8531 : _7593;
    assign _8533 = _7880 ? _7593 : _8532;
    assign _8534 = _7886 ? _7593 : _8533;
    assign _8535 = _7890 ? _7593 : _8534;
    assign _8536 = _7894 ? _7593 : _8535;
    assign _8537 = _7910 ? _7593 : _8536;
    assign _8538 = _7925 ? _7593 : _8537;
    assign _8539 = _6743 == _6738;
    assign _8540 = _8539 ? _8538 : _7593;
    assign _7591 = _8540;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7593 <= vdd;
        else
            _7593 <= _7591;
    end
    assign _7848 = _7839[8:8];
    assign _8521 = vdd ? _7848 : _7596;
    assign _8522 = _7874 ? _8521 : _7596;
    assign _8523 = _7880 ? _7596 : _8522;
    assign _8524 = _7886 ? _7596 : _8523;
    assign _8525 = _7890 ? _7596 : _8524;
    assign _8526 = _7894 ? _7596 : _8525;
    assign _8527 = _7910 ? _7596 : _8526;
    assign _8528 = _7925 ? _7596 : _8527;
    assign _8529 = _6743 == _6738;
    assign _8530 = _8529 ? _8528 : _7596;
    assign _7594 = _8530;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7596 <= vdd;
        else
            _7596 <= _7594;
    end
    assign _7849 = _7839[9:9];
    assign _8511 = vdd ? _7849 : _7599;
    assign _8512 = _7874 ? _8511 : _7599;
    assign _8513 = _7880 ? _7599 : _8512;
    assign _8514 = _7886 ? _7599 : _8513;
    assign _8515 = _7890 ? _7599 : _8514;
    assign _8516 = _7894 ? _7599 : _8515;
    assign _8517 = _7910 ? _7599 : _8516;
    assign _8518 = _7925 ? _7599 : _8517;
    assign _8519 = _6743 == _6738;
    assign _8520 = _8519 ? _8518 : _7599;
    assign _7597 = _8520;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7599 <= vdd;
        else
            _7599 <= _7597;
    end
    assign _7850 = _7839[10:10];
    assign _8501 = vdd ? _7850 : _7602;
    assign _8502 = _7874 ? _8501 : _7602;
    assign _8503 = _7880 ? _7602 : _8502;
    assign _8504 = _7886 ? _7602 : _8503;
    assign _8505 = _7890 ? _7602 : _8504;
    assign _8506 = _7894 ? _7602 : _8505;
    assign _8507 = _7910 ? _7602 : _8506;
    assign _8508 = _7925 ? _7602 : _8507;
    assign _8509 = _6743 == _6738;
    assign _8510 = _8509 ? _8508 : _7602;
    assign _7600 = _8510;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7602 <= vdd;
        else
            _7602 <= _7600;
    end
    assign _7851 = _7839[11:11];
    assign _8491 = vdd ? _7851 : _7605;
    assign _8492 = _7874 ? _8491 : _7605;
    assign _8493 = _7880 ? _7605 : _8492;
    assign _8494 = _7886 ? _7605 : _8493;
    assign _8495 = _7890 ? _7605 : _8494;
    assign _8496 = _7894 ? _7605 : _8495;
    assign _8497 = _7910 ? _7605 : _8496;
    assign _8498 = _7925 ? _7605 : _8497;
    assign _8499 = _6743 == _6738;
    assign _8500 = _8499 ? _8498 : _7605;
    assign _7603 = _8500;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7605 <= vdd;
        else
            _7605 <= _7603;
    end
    assign _7852 = _7839[12:12];
    assign _8481 = vdd ? _7852 : _7608;
    assign _8482 = _7874 ? _8481 : _7608;
    assign _8483 = _7880 ? _7608 : _8482;
    assign _8484 = _7886 ? _7608 : _8483;
    assign _8485 = _7890 ? _7608 : _8484;
    assign _8486 = _7894 ? _7608 : _8485;
    assign _8487 = _7910 ? _7608 : _8486;
    assign _8488 = _7925 ? _7608 : _8487;
    assign _8489 = _6743 == _6738;
    assign _8490 = _8489 ? _8488 : _7608;
    assign _7606 = _8490;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7608 <= vdd;
        else
            _7608 <= _7606;
    end
    assign _7853 = _7839[13:13];
    assign _8471 = vdd ? _7853 : _7611;
    assign _8472 = _7874 ? _8471 : _7611;
    assign _8473 = _7880 ? _7611 : _8472;
    assign _8474 = _7886 ? _7611 : _8473;
    assign _8475 = _7890 ? _7611 : _8474;
    assign _8476 = _7894 ? _7611 : _8475;
    assign _8477 = _7910 ? _7611 : _8476;
    assign _8478 = _7925 ? _7611 : _8477;
    assign _8479 = _6743 == _6738;
    assign _8480 = _8479 ? _8478 : _7611;
    assign _7609 = _8480;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7611 <= vdd;
        else
            _7611 <= _7609;
    end
    assign _7854 = _7839[14:14];
    assign _8461 = vdd ? _7854 : _7614;
    assign _8462 = _7874 ? _8461 : _7614;
    assign _8463 = _7880 ? _7614 : _8462;
    assign _8464 = _7886 ? _7614 : _8463;
    assign _8465 = _7890 ? _7614 : _8464;
    assign _8466 = _7894 ? _7614 : _8465;
    assign _8467 = _7910 ? _7614 : _8466;
    assign _8468 = _7925 ? _7614 : _8467;
    assign _8469 = _6743 == _6738;
    assign _8470 = _8469 ? _8468 : _7614;
    assign _7612 = _8470;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7614 <= vdd;
        else
            _7614 <= _7612;
    end
    assign _7855 = _7839[15:15];
    assign _8451 = vdd ? _7855 : _7617;
    assign _8452 = _7874 ? _8451 : _7617;
    assign _8453 = _7880 ? _7617 : _8452;
    assign _8454 = _7886 ? _7617 : _8453;
    assign _8455 = _7890 ? _7617 : _8454;
    assign _8456 = _7894 ? _7617 : _8455;
    assign _8457 = _7910 ? _7617 : _8456;
    assign _8458 = _7925 ? _7617 : _8457;
    assign _8459 = _6743 == _6738;
    assign _8460 = _8459 ? _8458 : _7617;
    assign _7615 = _8460;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7617 <= vdd;
        else
            _7617 <= _7615;
    end
    assign _7856 = _7839[16:16];
    assign _8441 = vdd ? _7856 : _7620;
    assign _8442 = _7874 ? _8441 : _7620;
    assign _8443 = _7880 ? _7620 : _8442;
    assign _8444 = _7886 ? _7620 : _8443;
    assign _8445 = _7890 ? _7620 : _8444;
    assign _8446 = _7894 ? _7620 : _8445;
    assign _8447 = _7910 ? _7620 : _8446;
    assign _8448 = _7925 ? _7620 : _8447;
    assign _8449 = _6743 == _6738;
    assign _8450 = _8449 ? _8448 : _7620;
    assign _7618 = _8450;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7620 <= vdd;
        else
            _7620 <= _7618;
    end
    assign _7857 = _7839[17:17];
    assign _8431 = vdd ? _7857 : _7623;
    assign _8432 = _7874 ? _8431 : _7623;
    assign _8433 = _7880 ? _7623 : _8432;
    assign _8434 = _7886 ? _7623 : _8433;
    assign _8435 = _7890 ? _7623 : _8434;
    assign _8436 = _7894 ? _7623 : _8435;
    assign _8437 = _7910 ? _7623 : _8436;
    assign _8438 = _7925 ? _7623 : _8437;
    assign _8439 = _6743 == _6738;
    assign _8440 = _8439 ? _8438 : _7623;
    assign _7621 = _8440;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7623 <= vdd;
        else
            _7623 <= _7621;
    end
    assign _7858 = _7839[18:18];
    assign _8421 = vdd ? _7858 : _7626;
    assign _8422 = _7874 ? _8421 : _7626;
    assign _8423 = _7880 ? _7626 : _8422;
    assign _8424 = _7886 ? _7626 : _8423;
    assign _8425 = _7890 ? _7626 : _8424;
    assign _8426 = _7894 ? _7626 : _8425;
    assign _8427 = _7910 ? _7626 : _8426;
    assign _8428 = _7925 ? _7626 : _8427;
    assign _8429 = _6743 == _6738;
    assign _8430 = _8429 ? _8428 : _7626;
    assign _7624 = _8430;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7626 <= vdd;
        else
            _7626 <= _7624;
    end
    assign _7859 = _7839[19:19];
    assign _8411 = vdd ? _7859 : _7629;
    assign _8412 = _7874 ? _8411 : _7629;
    assign _8413 = _7880 ? _7629 : _8412;
    assign _8414 = _7886 ? _7629 : _8413;
    assign _8415 = _7890 ? _7629 : _8414;
    assign _8416 = _7894 ? _7629 : _8415;
    assign _8417 = _7910 ? _7629 : _8416;
    assign _8418 = _7925 ? _7629 : _8417;
    assign _8419 = _6743 == _6738;
    assign _8420 = _8419 ? _8418 : _7629;
    assign _7627 = _8420;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7629 <= vdd;
        else
            _7629 <= _7627;
    end
    assign _7860 = _7839[20:20];
    assign _8401 = vdd ? _7860 : _7632;
    assign _8402 = _7874 ? _8401 : _7632;
    assign _8403 = _7880 ? _7632 : _8402;
    assign _8404 = _7886 ? _7632 : _8403;
    assign _8405 = _7890 ? _7632 : _8404;
    assign _8406 = _7894 ? _7632 : _8405;
    assign _8407 = _7910 ? _7632 : _8406;
    assign _8408 = _7925 ? _7632 : _8407;
    assign _8409 = _6743 == _6738;
    assign _8410 = _8409 ? _8408 : _7632;
    assign _7630 = _8410;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7632 <= vdd;
        else
            _7632 <= _7630;
    end
    assign _7861 = _7839[21:21];
    assign _8391 = vdd ? _7861 : _7635;
    assign _8392 = _7874 ? _8391 : _7635;
    assign _8393 = _7880 ? _7635 : _8392;
    assign _8394 = _7886 ? _7635 : _8393;
    assign _8395 = _7890 ? _7635 : _8394;
    assign _8396 = _7894 ? _7635 : _8395;
    assign _8397 = _7910 ? _7635 : _8396;
    assign _8398 = _7925 ? _7635 : _8397;
    assign _8399 = _6743 == _6738;
    assign _8400 = _8399 ? _8398 : _7635;
    assign _7633 = _8400;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7635 <= vdd;
        else
            _7635 <= _7633;
    end
    assign _7862 = _7839[22:22];
    assign _8381 = vdd ? _7862 : _7638;
    assign _8382 = _7874 ? _8381 : _7638;
    assign _8383 = _7880 ? _7638 : _8382;
    assign _8384 = _7886 ? _7638 : _8383;
    assign _8385 = _7890 ? _7638 : _8384;
    assign _8386 = _7894 ? _7638 : _8385;
    assign _8387 = _7910 ? _7638 : _8386;
    assign _8388 = _7925 ? _7638 : _8387;
    assign _8389 = _6743 == _6738;
    assign _8390 = _8389 ? _8388 : _7638;
    assign _7636 = _8390;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7638 <= vdd;
        else
            _7638 <= _7636;
    end
    assign _7863 = _7839[23:23];
    assign _8371 = vdd ? _7863 : _7641;
    assign _8372 = _7874 ? _8371 : _7641;
    assign _8373 = _7880 ? _7641 : _8372;
    assign _8374 = _7886 ? _7641 : _8373;
    assign _8375 = _7890 ? _7641 : _8374;
    assign _8376 = _7894 ? _7641 : _8375;
    assign _8377 = _7910 ? _7641 : _8376;
    assign _8378 = _7925 ? _7641 : _8377;
    assign _8379 = _6743 == _6738;
    assign _8380 = _8379 ? _8378 : _7641;
    assign _7639 = _8380;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7641 <= vdd;
        else
            _7641 <= _7639;
    end
    assign _7864 = _7839[24:24];
    assign _8361 = vdd ? _7864 : _7644;
    assign _8362 = _7874 ? _8361 : _7644;
    assign _8363 = _7880 ? _7644 : _8362;
    assign _8364 = _7886 ? _7644 : _8363;
    assign _8365 = _7890 ? _7644 : _8364;
    assign _8366 = _7894 ? _7644 : _8365;
    assign _8367 = _7910 ? _7644 : _8366;
    assign _8368 = _7925 ? _7644 : _8367;
    assign _8369 = _6743 == _6738;
    assign _8370 = _8369 ? _8368 : _7644;
    assign _7642 = _8370;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7644 <= vdd;
        else
            _7644 <= _7642;
    end
    assign _7865 = _7839[25:25];
    assign _8351 = vdd ? _7865 : _7647;
    assign _8352 = _7874 ? _8351 : _7647;
    assign _8353 = _7880 ? _7647 : _8352;
    assign _8354 = _7886 ? _7647 : _8353;
    assign _8355 = _7890 ? _7647 : _8354;
    assign _8356 = _7894 ? _7647 : _8355;
    assign _8357 = _7910 ? _7647 : _8356;
    assign _8358 = _7925 ? _7647 : _8357;
    assign _8359 = _6743 == _6738;
    assign _8360 = _8359 ? _8358 : _7647;
    assign _7645 = _8360;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7647 <= vdd;
        else
            _7647 <= _7645;
    end
    assign _7866 = _7839[26:26];
    assign _8341 = vdd ? _7866 : _7650;
    assign _8342 = _7874 ? _8341 : _7650;
    assign _8343 = _7880 ? _7650 : _8342;
    assign _8344 = _7886 ? _7650 : _8343;
    assign _8345 = _7890 ? _7650 : _8344;
    assign _8346 = _7894 ? _7650 : _8345;
    assign _8347 = _7910 ? _7650 : _8346;
    assign _8348 = _7925 ? _7650 : _8347;
    assign _8349 = _6743 == _6738;
    assign _8350 = _8349 ? _8348 : _7650;
    assign _7648 = _8350;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7650 <= vdd;
        else
            _7650 <= _7648;
    end
    assign _7867 = _7839[27:27];
    assign _8331 = vdd ? _7867 : _7653;
    assign _8332 = _7874 ? _8331 : _7653;
    assign _8333 = _7880 ? _7653 : _8332;
    assign _8334 = _7886 ? _7653 : _8333;
    assign _8335 = _7890 ? _7653 : _8334;
    assign _8336 = _7894 ? _7653 : _8335;
    assign _8337 = _7910 ? _7653 : _8336;
    assign _8338 = _7925 ? _7653 : _8337;
    assign _8339 = _6743 == _6738;
    assign _8340 = _8339 ? _8338 : _7653;
    assign _7651 = _8340;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7653 <= vdd;
        else
            _7653 <= _7651;
    end
    assign _7868 = _7839[28:28];
    assign _8321 = vdd ? _7868 : _7656;
    assign _8322 = _7874 ? _8321 : _7656;
    assign _8323 = _7880 ? _7656 : _8322;
    assign _8324 = _7886 ? _7656 : _8323;
    assign _8325 = _7890 ? _7656 : _8324;
    assign _8326 = _7894 ? _7656 : _8325;
    assign _8327 = _7910 ? _7656 : _8326;
    assign _8328 = _7925 ? _7656 : _8327;
    assign _8329 = _6743 == _6738;
    assign _8330 = _8329 ? _8328 : _7656;
    assign _7654 = _8330;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7656 <= vdd;
        else
            _7656 <= _7654;
    end
    assign _7869 = _7839[29:29];
    assign _8311 = vdd ? _7869 : _7659;
    assign _8312 = _7874 ? _8311 : _7659;
    assign _8313 = _7880 ? _7659 : _8312;
    assign _8314 = _7886 ? _7659 : _8313;
    assign _8315 = _7890 ? _7659 : _8314;
    assign _8316 = _7894 ? _7659 : _8315;
    assign _8317 = _7910 ? _7659 : _8316;
    assign _8318 = _7925 ? _7659 : _8317;
    assign _8319 = _6743 == _6738;
    assign _8320 = _8319 ? _8318 : _7659;
    assign _7657 = _8320;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7659 <= vdd;
        else
            _7659 <= _7657;
    end
    assign _7870 = _7839[30:30];
    assign _8301 = vdd ? _7870 : _7662;
    assign _8302 = _7874 ? _8301 : _7662;
    assign _8303 = _7880 ? _7662 : _8302;
    assign _8304 = _7886 ? _7662 : _8303;
    assign _8305 = _7890 ? _7662 : _8304;
    assign _8306 = _7894 ? _7662 : _8305;
    assign _8307 = _7910 ? _7662 : _8306;
    assign _8308 = _7925 ? _7662 : _8307;
    assign _8309 = _6743 == _6738;
    assign _8310 = _8309 ? _8308 : _7662;
    assign _7660 = _8310;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7662 <= vdd;
        else
            _7662 <= _7660;
    end
    assign _7871 = _7839[31:31];
    assign _8291 = vdd ? _7871 : _7665;
    assign _8292 = _7874 ? _8291 : _7665;
    assign _8293 = _7880 ? _7665 : _8292;
    assign _8294 = _7886 ? _7665 : _8293;
    assign _8295 = _7890 ? _7665 : _8294;
    assign _8296 = _7894 ? _7665 : _8295;
    assign _8297 = _7910 ? _7665 : _8296;
    assign _8298 = _7925 ? _7665 : _8297;
    assign _8299 = _6743 == _6738;
    assign _8300 = _8299 ? _8298 : _7665;
    assign _7663 = _8300;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7665 <= vdd;
        else
            _7665 <= _7663;
    end
    assign _7666 = { _7665, _7662, _7659, _7656, _7653, _7650, _7647, _7644, _7641, _7638, _7635, _7632, _7629, _7626, _7623, _7620, _7617, _7614, _7611, _7608, _7605, _7602, _7599, _7596, _7593, _7590, _7587, _7584, _7581, _7578, _7575, _7572 };
    assign _7796 = _7569 & _7666;
    assign _8660 = _7802 ? _7796 : _7569;
    assign _8661 = _7806 ? _7569 : _8660;
    assign _8662 = _7492 ? _7569 : _8661;
    assign _8663 = _7484 ? _7569 : _8662;
    assign _8088 = _7673 - _8087;
    assign _8090 = _8088 == _8089;
    assign _8658 = _8090 ? _8086 : _8657;
    assign _8105 = irq[0:0];
    assign _8106 = _38[0:0];
    assign _8107 = _7536[0:0];
    assign _8108 = _8107 & _8106;
    assign _8109 = _8108 | _8105;
    assign _8657 = vdd ? _8109 : gnd;
    assign _8269 = _7838 ? _7820 : _8268;
    assign _8270 = _7874 ? _8268 : _8269;
    assign _8271 = _7880 ? _8268 : _8270;
    assign _8272 = _7886 ? _8268 : _8271;
    assign _8273 = _7890 ? _8268 : _8272;
    assign _8274 = _7894 ? _8268 : _8273;
    assign _8275 = _7910 ? _8268 : _8274;
    assign _8276 = _7925 ? _8268 : _8275;
    assign _8085 = _7673 - _8084;
    assign _8268 = _8095 ? _8085 : _7673;
    assign _8277 = _6743 == _6738;
    assign _8278 = _8277 ? _8276 : _8268;
    assign _7671 = _8278;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7673 <= _7670;
        else
            _7673 <= _7671;
    end
    assign _8092 = _7673 == _8091;
    assign _8093 = ~ _8092;
    assign _8094 = vdd & vdd;
    assign _8095 = _8094 & _8093;
    assign _8659 = _8095 ? _8658 : _8657;
    assign _7537 = _8659;
    assign _7917 = ~ _7532;
    assign _7918 = ~ _7575;
    assign _7919 = vdd & _7918;
    assign _7920 = _7919 & _7917;
    assign _8642 = _7920 ? _7916 : _8641;
    assign _8643 = _7464 ? _8642 : _8641;
    assign _8644 = _5634 ? _8641 : _8643;
    assign _8645 = vdd ? _8644 : _8641;
    assign _7912 = ~ _7532;
    assign _7913 = ~ _7575;
    assign _7914 = vdd & _7913;
    assign _7915 = _7914 & _7912;
    assign _8646 = _7915 ? _7911 : _8641;
    assign _8647 = vdd ? _8645 : _8646;
    assign _8648 = _7925 ? _8647 : _8641;
    assign _7932 = ~ _7532;
    assign _7376 = _7200[35:35];
    assign _7377 = _6810 & _7376;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7380 <= _7378;
        else
            if (_7377)
                _7380 <= _6809;
    end
    assign _7371 = _7200[34:34];
    assign _7372 = _6810 & _7371;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7375 <= _7373;
        else
            if (_7372)
                _7375 <= _6809;
    end
    assign _7366 = _7200[33:33];
    assign _7367 = _6810 & _7366;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7370 <= _7368;
        else
            if (_7367)
                _7370 <= _6809;
    end
    assign _7361 = _7200[32:32];
    assign _7362 = _6810 & _7361;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7365 <= _7363;
        else
            if (_7362)
                _7365 <= _6809;
    end
    assign _7356 = _7200[31:31];
    assign _7357 = _6810 & _7356;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7360 <= _7358;
        else
            if (_7357)
                _7360 <= _6809;
    end
    assign _7351 = _7200[30:30];
    assign _7352 = _6810 & _7351;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7355 <= _7353;
        else
            if (_7352)
                _7355 <= _6809;
    end
    assign _7346 = _7200[29:29];
    assign _7347 = _6810 & _7346;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7350 <= _7348;
        else
            if (_7347)
                _7350 <= _6809;
    end
    assign _7341 = _7200[28:28];
    assign _7342 = _6810 & _7341;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7345 <= _7343;
        else
            if (_7342)
                _7345 <= _6809;
    end
    assign _7336 = _7200[27:27];
    assign _7337 = _6810 & _7336;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7340 <= _7338;
        else
            if (_7337)
                _7340 <= _6809;
    end
    assign _7331 = _7200[26:26];
    assign _7332 = _6810 & _7331;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7335 <= _7333;
        else
            if (_7332)
                _7335 <= _6809;
    end
    assign _7326 = _7200[25:25];
    assign _7327 = _6810 & _7326;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7330 <= _7328;
        else
            if (_7327)
                _7330 <= _6809;
    end
    assign _7321 = _7200[24:24];
    assign _7322 = _6810 & _7321;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7325 <= _7323;
        else
            if (_7322)
                _7325 <= _6809;
    end
    assign _7316 = _7200[23:23];
    assign _7317 = _6810 & _7316;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7320 <= _7318;
        else
            if (_7317)
                _7320 <= _6809;
    end
    assign _7311 = _7200[22:22];
    assign _7312 = _6810 & _7311;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7315 <= _7313;
        else
            if (_7312)
                _7315 <= _6809;
    end
    assign _7306 = _7200[21:21];
    assign _7307 = _6810 & _7306;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7310 <= _7308;
        else
            if (_7307)
                _7310 <= _6809;
    end
    assign _7301 = _7200[20:20];
    assign _7302 = _6810 & _7301;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7305 <= _7303;
        else
            if (_7302)
                _7305 <= _6809;
    end
    assign _7296 = _7200[19:19];
    assign _7297 = _6810 & _7296;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7300 <= _7298;
        else
            if (_7297)
                _7300 <= _6809;
    end
    assign _7291 = _7200[18:18];
    assign _7292 = _6810 & _7291;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7295 <= _7293;
        else
            if (_7292)
                _7295 <= _6809;
    end
    assign _7286 = _7200[17:17];
    assign _7287 = _6810 & _7286;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7290 <= _7288;
        else
            if (_7287)
                _7290 <= _6809;
    end
    assign _7281 = _7200[16:16];
    assign _7282 = _6810 & _7281;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7285 <= _7283;
        else
            if (_7282)
                _7285 <= _6809;
    end
    assign _7276 = _7200[15:15];
    assign _7277 = _6810 & _7276;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7280 <= _7278;
        else
            if (_7277)
                _7280 <= _6809;
    end
    assign _7271 = _7200[14:14];
    assign _7272 = _6810 & _7271;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7275 <= _7273;
        else
            if (_7272)
                _7275 <= _6809;
    end
    assign _7266 = _7200[13:13];
    assign _7267 = _6810 & _7266;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7270 <= _7268;
        else
            if (_7267)
                _7270 <= _6809;
    end
    assign _7261 = _7200[12:12];
    assign _7262 = _6810 & _7261;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7265 <= _7263;
        else
            if (_7262)
                _7265 <= _6809;
    end
    assign _7256 = _7200[11:11];
    assign _7257 = _6810 & _7256;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7260 <= _7258;
        else
            if (_7257)
                _7260 <= _6809;
    end
    assign _7251 = _7200[10:10];
    assign _7252 = _6810 & _7251;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7255 <= _7253;
        else
            if (_7252)
                _7255 <= _6809;
    end
    assign _7246 = _7200[9:9];
    assign _7247 = _6810 & _7246;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7250 <= _7248;
        else
            if (_7247)
                _7250 <= _6809;
    end
    assign _7241 = _7200[8:8];
    assign _7242 = _6810 & _7241;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7245 <= _7243;
        else
            if (_7242)
                _7245 <= _6809;
    end
    assign _7236 = _7200[7:7];
    assign _7237 = _6810 & _7236;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7240 <= _7238;
        else
            if (_7237)
                _7240 <= _6809;
    end
    assign _7231 = _7200[6:6];
    assign _7232 = _6810 & _7231;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7235 <= _7233;
        else
            if (_7232)
                _7235 <= _6809;
    end
    assign _7226 = _7200[5:5];
    assign _7227 = _6810 & _7226;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7230 <= _7228;
        else
            if (_7227)
                _7230 <= _6809;
    end
    assign _7221 = _7200[4:4];
    assign _7222 = _6810 & _7221;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7225 <= _7223;
        else
            if (_7222)
                _7225 <= _6809;
    end
    assign _7216 = _7200[3:3];
    assign _7217 = _6810 & _7216;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7220 <= _7218;
        else
            if (_7217)
                _7220 <= _6809;
    end
    assign _7211 = _7200[2:2];
    assign _7212 = _6810 & _7211;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7215 <= _7213;
        else
            if (_7212)
                _7215 <= _6809;
    end
    assign _6817 = ~ _6811;
    assign _6820 = _6818 & _6817;
    assign _6828 = _6824 & _6820;
    assign _6848 = _6840 & _6828;
    assign _6896 = _6880 & _6848;
    assign _7008 = _6976 & _6896;
    assign _6818 = ~ _6812;
    assign _6819 = _6818 & _6811;
    assign _6827 = _6824 & _6819;
    assign _6847 = _6840 & _6827;
    assign _6895 = _6880 & _6847;
    assign _7007 = _6976 & _6895;
    assign _6821 = ~ _6811;
    assign _6823 = _6812 & _6821;
    assign _6826 = _6824 & _6823;
    assign _6846 = _6840 & _6826;
    assign _6894 = _6880 & _6846;
    assign _7006 = _6976 & _6894;
    assign _6822 = _6812 & _6811;
    assign _6824 = ~ _6813;
    assign _6825 = _6824 & _6822;
    assign _6845 = _6840 & _6825;
    assign _6893 = _6880 & _6845;
    assign _7005 = _6976 & _6893;
    assign _6829 = ~ _6811;
    assign _6832 = _6830 & _6829;
    assign _6839 = _6813 & _6832;
    assign _6844 = _6840 & _6839;
    assign _6892 = _6880 & _6844;
    assign _7004 = _6976 & _6892;
    assign _6830 = ~ _6812;
    assign _6831 = _6830 & _6811;
    assign _6838 = _6813 & _6831;
    assign _6843 = _6840 & _6838;
    assign _6891 = _6880 & _6843;
    assign _7003 = _6976 & _6891;
    assign _6833 = ~ _6811;
    assign _6835 = _6812 & _6833;
    assign _6837 = _6813 & _6835;
    assign _6842 = _6840 & _6837;
    assign _6890 = _6880 & _6842;
    assign _7002 = _6976 & _6890;
    assign _6834 = _6812 & _6811;
    assign _6836 = _6813 & _6834;
    assign _6840 = ~ _6814;
    assign _6841 = _6840 & _6836;
    assign _6889 = _6880 & _6841;
    assign _7001 = _6976 & _6889;
    assign _6849 = ~ _6811;
    assign _6852 = _6850 & _6849;
    assign _6860 = _6856 & _6852;
    assign _6879 = _6814 & _6860;
    assign _6888 = _6880 & _6879;
    assign _7000 = _6976 & _6888;
    assign _6850 = ~ _6812;
    assign _6851 = _6850 & _6811;
    assign _6859 = _6856 & _6851;
    assign _6878 = _6814 & _6859;
    assign _6887 = _6880 & _6878;
    assign _6999 = _6976 & _6887;
    assign _6853 = ~ _6811;
    assign _6855 = _6812 & _6853;
    assign _6858 = _6856 & _6855;
    assign _6877 = _6814 & _6858;
    assign _6886 = _6880 & _6877;
    assign _6998 = _6976 & _6886;
    assign _6854 = _6812 & _6811;
    assign _6856 = ~ _6813;
    assign _6857 = _6856 & _6854;
    assign _6876 = _6814 & _6857;
    assign _6885 = _6880 & _6876;
    assign _6997 = _6976 & _6885;
    assign _6861 = ~ _6811;
    assign _6864 = _6862 & _6861;
    assign _6871 = _6813 & _6864;
    assign _6875 = _6814 & _6871;
    assign _6884 = _6880 & _6875;
    assign _6996 = _6976 & _6884;
    assign _6862 = ~ _6812;
    assign _6863 = _6862 & _6811;
    assign _6870 = _6813 & _6863;
    assign _6874 = _6814 & _6870;
    assign _6883 = _6880 & _6874;
    assign _6995 = _6976 & _6883;
    assign _6865 = ~ _6811;
    assign _6867 = _6812 & _6865;
    assign _6869 = _6813 & _6867;
    assign _6873 = _6814 & _6869;
    assign _6882 = _6880 & _6873;
    assign _6994 = _6976 & _6882;
    assign _6866 = _6812 & _6811;
    assign _6868 = _6813 & _6866;
    assign _6872 = _6814 & _6868;
    assign _6880 = ~ _6815;
    assign _6881 = _6880 & _6872;
    assign _6993 = _6976 & _6881;
    assign _6897 = ~ _6811;
    assign _6900 = _6898 & _6897;
    assign _6908 = _6904 & _6900;
    assign _6928 = _6920 & _6908;
    assign _6975 = _6815 & _6928;
    assign _6992 = _6976 & _6975;
    assign _6898 = ~ _6812;
    assign _6899 = _6898 & _6811;
    assign _6907 = _6904 & _6899;
    assign _6927 = _6920 & _6907;
    assign _6974 = _6815 & _6927;
    assign _6991 = _6976 & _6974;
    assign _6901 = ~ _6811;
    assign _6903 = _6812 & _6901;
    assign _6906 = _6904 & _6903;
    assign _6926 = _6920 & _6906;
    assign _6973 = _6815 & _6926;
    assign _6990 = _6976 & _6973;
    assign _6902 = _6812 & _6811;
    assign _6904 = ~ _6813;
    assign _6905 = _6904 & _6902;
    assign _6925 = _6920 & _6905;
    assign _6972 = _6815 & _6925;
    assign _6989 = _6976 & _6972;
    assign _6909 = ~ _6811;
    assign _6912 = _6910 & _6909;
    assign _6919 = _6813 & _6912;
    assign _6924 = _6920 & _6919;
    assign _6971 = _6815 & _6924;
    assign _6988 = _6976 & _6971;
    assign _6910 = ~ _6812;
    assign _6911 = _6910 & _6811;
    assign _6918 = _6813 & _6911;
    assign _6923 = _6920 & _6918;
    assign _6970 = _6815 & _6923;
    assign _6987 = _6976 & _6970;
    assign _6913 = ~ _6811;
    assign _6915 = _6812 & _6913;
    assign _6917 = _6813 & _6915;
    assign _6922 = _6920 & _6917;
    assign _6969 = _6815 & _6922;
    assign _6986 = _6976 & _6969;
    assign _6914 = _6812 & _6811;
    assign _6916 = _6813 & _6914;
    assign _6920 = ~ _6814;
    assign _6921 = _6920 & _6916;
    assign _6968 = _6815 & _6921;
    assign _6985 = _6976 & _6968;
    assign _6929 = ~ _6811;
    assign _6932 = _6930 & _6929;
    assign _6940 = _6936 & _6932;
    assign _6959 = _6814 & _6940;
    assign _6967 = _6815 & _6959;
    assign _6984 = _6976 & _6967;
    assign _6930 = ~ _6812;
    assign _6931 = _6930 & _6811;
    assign _6939 = _6936 & _6931;
    assign _6958 = _6814 & _6939;
    assign _6966 = _6815 & _6958;
    assign _6983 = _6976 & _6966;
    assign _6933 = ~ _6811;
    assign _6935 = _6812 & _6933;
    assign _6938 = _6936 & _6935;
    assign _6957 = _6814 & _6938;
    assign _6965 = _6815 & _6957;
    assign _6982 = _6976 & _6965;
    assign _6934 = _6812 & _6811;
    assign _6936 = ~ _6813;
    assign _6937 = _6936 & _6934;
    assign _6956 = _6814 & _6937;
    assign _6964 = _6815 & _6956;
    assign _6981 = _6976 & _6964;
    assign _6941 = ~ _6811;
    assign _6944 = _6942 & _6941;
    assign _6951 = _6813 & _6944;
    assign _6955 = _6814 & _6951;
    assign _6963 = _6815 & _6955;
    assign _6980 = _6976 & _6963;
    assign _6942 = ~ _6812;
    assign _6943 = _6942 & _6811;
    assign _6950 = _6813 & _6943;
    assign _6954 = _6814 & _6950;
    assign _6962 = _6815 & _6954;
    assign _6979 = _6976 & _6962;
    assign _6945 = ~ _6811;
    assign _6947 = _6812 & _6945;
    assign _6949 = _6813 & _6947;
    assign _6953 = _6814 & _6949;
    assign _6961 = _6815 & _6953;
    assign _6978 = _6976 & _6961;
    assign _6946 = _6812 & _6811;
    assign _6948 = _6813 & _6946;
    assign _6952 = _6814 & _6948;
    assign _6960 = _6815 & _6952;
    assign _6976 = ~ _6816;
    assign _6977 = _6976 & _6960;
    assign _7009 = ~ _6811;
    assign _7012 = _7010 & _7009;
    assign _7020 = _7016 & _7012;
    assign _7040 = _7032 & _7020;
    assign _7088 = _7072 & _7040;
    assign _7199 = _6816 & _7088;
    assign _7010 = ~ _6812;
    assign _7011 = _7010 & _6811;
    assign _7019 = _7016 & _7011;
    assign _7039 = _7032 & _7019;
    assign _7087 = _7072 & _7039;
    assign _7198 = _6816 & _7087;
    assign _7013 = ~ _6811;
    assign _7015 = _6812 & _7013;
    assign _7018 = _7016 & _7015;
    assign _7038 = _7032 & _7018;
    assign _7086 = _7072 & _7038;
    assign _7197 = _6816 & _7086;
    assign _7014 = _6812 & _6811;
    assign _7016 = ~ _6813;
    assign _7017 = _7016 & _7014;
    assign _7037 = _7032 & _7017;
    assign _7085 = _7072 & _7037;
    assign _7196 = _6816 & _7085;
    assign _7021 = ~ _6811;
    assign _7024 = _7022 & _7021;
    assign _7031 = _6813 & _7024;
    assign _7036 = _7032 & _7031;
    assign _7084 = _7072 & _7036;
    assign _7195 = _6816 & _7084;
    assign _7022 = ~ _6812;
    assign _7023 = _7022 & _6811;
    assign _7030 = _6813 & _7023;
    assign _7035 = _7032 & _7030;
    assign _7083 = _7072 & _7035;
    assign _7194 = _6816 & _7083;
    assign _7025 = ~ _6811;
    assign _7027 = _6812 & _7025;
    assign _7029 = _6813 & _7027;
    assign _7034 = _7032 & _7029;
    assign _7082 = _7072 & _7034;
    assign _7193 = _6816 & _7082;
    assign _7026 = _6812 & _6811;
    assign _7028 = _6813 & _7026;
    assign _7032 = ~ _6814;
    assign _7033 = _7032 & _7028;
    assign _7081 = _7072 & _7033;
    assign _7192 = _6816 & _7081;
    assign _7041 = ~ _6811;
    assign _7044 = _7042 & _7041;
    assign _7052 = _7048 & _7044;
    assign _7071 = _6814 & _7052;
    assign _7080 = _7072 & _7071;
    assign _7191 = _6816 & _7080;
    assign _7042 = ~ _6812;
    assign _7043 = _7042 & _6811;
    assign _7051 = _7048 & _7043;
    assign _7070 = _6814 & _7051;
    assign _7079 = _7072 & _7070;
    assign _7190 = _6816 & _7079;
    assign _7045 = ~ _6811;
    assign _7047 = _6812 & _7045;
    assign _7050 = _7048 & _7047;
    assign _7069 = _6814 & _7050;
    assign _7078 = _7072 & _7069;
    assign _7189 = _6816 & _7078;
    assign _7046 = _6812 & _6811;
    assign _7048 = ~ _6813;
    assign _7049 = _7048 & _7046;
    assign _7068 = _6814 & _7049;
    assign _7077 = _7072 & _7068;
    assign _7188 = _6816 & _7077;
    assign _7053 = ~ _6811;
    assign _7056 = _7054 & _7053;
    assign _7063 = _6813 & _7056;
    assign _7067 = _6814 & _7063;
    assign _7076 = _7072 & _7067;
    assign _7187 = _6816 & _7076;
    assign _7054 = ~ _6812;
    assign _7055 = _7054 & _6811;
    assign _7062 = _6813 & _7055;
    assign _7066 = _6814 & _7062;
    assign _7075 = _7072 & _7066;
    assign _7186 = _6816 & _7075;
    assign _7057 = ~ _6811;
    assign _7059 = _6812 & _7057;
    assign _7061 = _6813 & _7059;
    assign _7065 = _6814 & _7061;
    assign _7074 = _7072 & _7065;
    assign _7185 = _6816 & _7074;
    assign _7058 = _6812 & _6811;
    assign _7060 = _6813 & _7058;
    assign _7064 = _6814 & _7060;
    assign _7072 = ~ _6815;
    assign _7073 = _7072 & _7064;
    assign _7184 = _6816 & _7073;
    assign _7089 = ~ _6811;
    assign _7092 = _7090 & _7089;
    assign _7100 = _7096 & _7092;
    assign _7120 = _7112 & _7100;
    assign _7167 = _6815 & _7120;
    assign _7183 = _6816 & _7167;
    assign _7090 = ~ _6812;
    assign _7091 = _7090 & _6811;
    assign _7099 = _7096 & _7091;
    assign _7119 = _7112 & _7099;
    assign _7166 = _6815 & _7119;
    assign _7182 = _6816 & _7166;
    assign _7093 = ~ _6811;
    assign _7095 = _6812 & _7093;
    assign _7098 = _7096 & _7095;
    assign _7118 = _7112 & _7098;
    assign _7165 = _6815 & _7118;
    assign _7181 = _6816 & _7165;
    assign _7094 = _6812 & _6811;
    assign _7096 = ~ _6813;
    assign _7097 = _7096 & _7094;
    assign _7117 = _7112 & _7097;
    assign _7164 = _6815 & _7117;
    assign _7180 = _6816 & _7164;
    assign _7101 = ~ _6811;
    assign _7104 = _7102 & _7101;
    assign _7111 = _6813 & _7104;
    assign _7116 = _7112 & _7111;
    assign _7163 = _6815 & _7116;
    assign _7179 = _6816 & _7163;
    assign _7102 = ~ _6812;
    assign _7103 = _7102 & _6811;
    assign _7110 = _6813 & _7103;
    assign _7115 = _7112 & _7110;
    assign _7162 = _6815 & _7115;
    assign _7178 = _6816 & _7162;
    assign _7105 = ~ _6811;
    assign _7107 = _6812 & _7105;
    assign _7109 = _6813 & _7107;
    assign _7114 = _7112 & _7109;
    assign _7161 = _6815 & _7114;
    assign _7177 = _6816 & _7161;
    assign _7106 = _6812 & _6811;
    assign _7108 = _6813 & _7106;
    assign _7112 = ~ _6814;
    assign _7113 = _7112 & _7108;
    assign _7160 = _6815 & _7113;
    assign _7176 = _6816 & _7160;
    assign _7121 = ~ _6811;
    assign _7124 = _7122 & _7121;
    assign _7132 = _7128 & _7124;
    assign _7151 = _6814 & _7132;
    assign _7159 = _6815 & _7151;
    assign _7175 = _6816 & _7159;
    assign _7122 = ~ _6812;
    assign _7123 = _7122 & _6811;
    assign _7131 = _7128 & _7123;
    assign _7150 = _6814 & _7131;
    assign _7158 = _6815 & _7150;
    assign _7174 = _6816 & _7158;
    assign _7125 = ~ _6811;
    assign _7127 = _6812 & _7125;
    assign _7130 = _7128 & _7127;
    assign _7149 = _6814 & _7130;
    assign _7157 = _6815 & _7149;
    assign _7173 = _6816 & _7157;
    assign _7126 = _6812 & _6811;
    assign _7128 = ~ _6813;
    assign _7129 = _7128 & _7126;
    assign _7148 = _6814 & _7129;
    assign _7156 = _6815 & _7148;
    assign _7172 = _6816 & _7156;
    assign _7133 = ~ _6811;
    assign _7136 = _7134 & _7133;
    assign _7143 = _6813 & _7136;
    assign _7147 = _6814 & _7143;
    assign _7155 = _6815 & _7147;
    assign _7171 = _6816 & _7155;
    assign _7134 = ~ _6812;
    assign _7135 = _7134 & _6811;
    assign _7142 = _6813 & _7135;
    assign _7146 = _6814 & _7142;
    assign _7154 = _6815 & _7146;
    assign _7170 = _6816 & _7154;
    assign _7137 = ~ _6811;
    assign _7139 = _6812 & _7137;
    assign _7141 = _6813 & _7139;
    assign _7145 = _6814 & _7141;
    assign _7153 = _6815 & _7145;
    assign _7169 = _6816 & _7153;
    assign _6811 = _6807[0:0];
    assign _6812 = _6807[1:1];
    assign _7138 = _6812 & _6811;
    assign _6813 = _6807[2:2];
    assign _7140 = _6813 & _7138;
    assign _6814 = _6807[3:3];
    assign _7144 = _6814 & _7140;
    assign _6815 = _6807[4:4];
    assign _7152 = _6815 & _7144;
    assign _7700 = _7528[0:0];
    assign _7705 = { _7703, _7700 };
    assign _7707 = _7706 | _7705;
    assign _7699 = _7528[0:0];
    assign _9113 = _7699 ? _7698 : _7697;
    assign _9114 = vdd ? _7707 : _9113;
    assign _6555 = _5653[11:7];
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6558 <= _6556;
        else
            if (_5841)
                _6558 <= _6555;
    end
    assign _6559 = { gnd, _6558 };
    assign _5642 = _6559;
    assign _9115 = _7789 ? _9114 : _5642;
    assign _7883 = _6807 | _7882;
    assign _9116 = _7886 ? _7883 : _6807;
    assign _9117 = _7890 ? _6807 : _9116;
    assign _9118 = _7894 ? _6807 : _9117;
    assign _9119 = _7910 ? _6807 : _9118;
    assign _9120 = _7925 ? _6807 : _9119;
    assign _9121 = _7948 ? _7947 : _6807;
    assign _9122 = _6743 == _6736;
    assign _9123 = _9122 ? _9121 : _6807;
    assign _9124 = _6743 == _6738;
    assign _9125 = _9124 ? _9120 : _9123;
    assign _9126 = _6743 == _6740;
    assign _9127 = _9126 ? _9115 : _9125;
    assign _6805 = _9127;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6807 <= _6804;
        else
            _6807 <= _6805;
    end
    assign _6816 = _6807[5:5];
    assign _7168 = _6816 & _7152;
    assign _7200 = { _7168, _7169, _7170, _7171, _7172, _7173, _7174, _7175, _7176, _7177, _7178, _7179, _7180, _7181, _7182, _7183, _7184, _7185, _7186, _7187, _7188, _7189, _7190, _7191, _7192, _7193, _7194, _7195, _7196, _7197, _7198, _7199, _6977, _6978, _6979, _6980, _6981, _6982, _6983, _6984, _6985, _6986, _6987, _6988, _6989, _6990, _6991, _6992, _6993, _6994, _6995, _6996, _6997, _6998, _6999, _7000, _7001, _7002, _7003, _7004, _7005, _7006, _7007, _7008 };
    assign _7206 = _7200[1:1];
    assign _9093 = vdd ? vdd : gnd;
    assign _9094 = vdd ? vdd : gnd;
    assign _9095 = vdd ? vdd : gnd;
    assign _9096 = vdd ? vdd : gnd;
    assign _7801 = _7528[1:1];
    assign _7802 = vdd & _7801;
    assign _9097 = _7802 ? _9096 : gnd;
    assign _7711 = _7528 == _7710;
    assign _7712 = _7711 ? _7709 : _7708;
    assign _7715 = _7528 == _7714;
    assign _7716 = _7715 ? _7713 : _7712;
    assign _8679 = _7789 ? _7716 : _7528;
    assign _8680 = _6743 == _6740;
    assign _8681 = _8680 ? _8679 : _7528;
    assign _7526 = _8681;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7528 <= _7525;
        else
            _7528 <= _7526;
    end
    assign _7805 = _7528[0:0];
    assign _7806 = vdd & _7805;
    assign _9098 = _7806 ? _9095 : _9097;
    assign _9099 = _7492 ? _9094 : _9098;
    assign _9100 = _7484 ? _9093 : _9099;
    assign _9101 = _6743 == _6740;
    assign _9102 = _9101 ? _9100 : gnd;
    assign _6810 = _9102;
    assign _7207 = _6810 & _7206;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7210 <= _7208;
        else
            if (_7207)
                _7210 <= _6809;
    end
    always @* begin
        case (_5641)
        0: _7382 <= _7205;
        1: _7382 <= _7210;
        2: _7382 <= _7215;
        3: _7382 <= _7220;
        4: _7382 <= _7225;
        5: _7382 <= _7230;
        6: _7382 <= _7235;
        7: _7382 <= _7240;
        8: _7382 <= _7245;
        9: _7382 <= _7250;
        10: _7382 <= _7255;
        11: _7382 <= _7260;
        12: _7382 <= _7265;
        13: _7382 <= _7270;
        14: _7382 <= _7275;
        15: _7382 <= _7280;
        16: _7382 <= _7285;
        17: _7382 <= _7290;
        18: _7382 <= _7295;
        19: _7382 <= _7300;
        20: _7382 <= _7305;
        21: _7382 <= _7310;
        22: _7382 <= _7315;
        23: _7382 <= _7320;
        24: _7382 <= _7325;
        25: _7382 <= _7330;
        26: _7382 <= _7335;
        27: _7382 <= _7340;
        28: _7382 <= _7345;
        29: _7382 <= _7350;
        30: _7382 <= _7355;
        31: _7382 <= _7360;
        32: _7382 <= _7365;
        33: _7382 <= _7370;
        34: _7382 <= _7375;
        default: _7382 <= _7380;
        endcase
    end
    assign _6466 = cx[4:0];
    assign _6467 = { vdd, _6466 };
    assign _6464 = _5653[19:15];
    assign cx = { gnd, _6464 };
    assign _6447 = _5653[31:25];
    assign _6449 = _6447 == _6448;
    assign _6450 = _5653[6:0];
    assign _6452 = _6450 == _6451;
    assign _6453 = _6452 & _6449;
    assign _6454 = _6453 & vdd;
    assign c0 = _6454 & vdd;
    assign _6468 = c0 ? _6467 : cx;
    assign _6456 = _5653[31:25];
    assign _6458 = _6456 == _6457;
    assign _6459 = _5653[6:0];
    assign _6461 = _6459 == _6460;
    assign _6462 = _6461 & _6458;
    assign c1 = _6462 & vdd;
    assign _6470 = c1 ? _6469 : _6468;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6554 <= _6552;
        else
            if (_5841)
                _6554 <= _6470;
    end
    assign _5641 = _6554;
    assign _7818 = _5641 == _7817;
    assign _7819 = ~ _7818;
    assign _7820 = _7819 ? _7382 : _7816;
    assign _7839 = _7820 | _37;
    assign _7841 = _7839[1:1];
    assign _8591 = vdd ? _7841 : _7575;
    assign _8592 = _7874 ? _8591 : _7575;
    assign _8593 = _7880 ? _7575 : _8592;
    assign _8594 = _7886 ? _7575 : _8593;
    assign _8595 = _7890 ? _7575 : _8594;
    assign _8596 = _7894 ? _7575 : _8595;
    assign _8597 = _7910 ? _7575 : _8596;
    assign _8598 = _7925 ? _7575 : _8597;
    assign _8599 = _6743 == _6738;
    assign _8600 = _8599 ? _8598 : _7575;
    assign _7573 = _8600;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7575 <= vdd;
        else
            _7575 <= _7573;
    end
    assign _7933 = ~ _7575;
    assign _7934 = vdd & _7933;
    assign _7935 = _7934 & _7932;
    assign _8649 = _7935 ? _7931 : _8641;
    assign _8102 = _7468 - _8101;
    assign _9082 = _7468[0:0];
    assign _9083 = _7468[1:1];
    assign _9084 = _7468[2:2];
    assign _9085 = _7468[3:3];
    assign _9086 = _9085 | _9084;
    assign _9087 = _9086 | _9083;
    assign _9088 = _9087 | _9082;
    assign _9089 = _9088 ? _8102 : _7468;
    assign _5830 = vdd & _5719;
    assign _5831 = gnd & pcpi_wait;
    assign _5832 = _5831 | _5830;
    assign _5635 = _5832;
    assign _8103 = ~ _5635;
    assign _8104 = _6767 & _8103;
    assign _9090 = _8104 ? _9089 : _8100;
    assign _9091 = vdd ? _9090 : _7468;
    assign _7466 = _9091;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7468 <= _7465;
        else
            _7468 <= _7466;
    end
    assign _8099 = _7468 == _8098;
    assign _9092 = vdd ? _8099 : _7464;
    assign _7462 = _9092;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7464 <= _7461;
        else
            _7464 <= _7462;
    end
    assign _8650 = _7464 ? _8649 : _8641;
    assign _8651 = _5634 ? _8641 : _8650;
    assign _8652 = _7940 ? _8651 : _8641;
    assign _8110 = irq[1:1];
    assign _8111 = _38[1:1];
    assign _8112 = _7536[1:1];
    assign _8113 = _8112 & _8111;
    assign _8114 = _8113 | _8110;
    assign _8641 = vdd ? _8114 : gnd;
    assign _8653 = _6743 == _6737;
    assign _8654 = _8653 ? _8652 : _8641;
    assign _8655 = _6743 == _6738;
    assign _8656 = _8655 ? _8648 : _8654;
    assign _7538 = _8656;
    assign _8115 = irq[2:2];
    assign _8116 = _38[2:2];
    assign _8117 = _7536[2:2];
    assign _8118 = _8117 & _8116;
    assign _8119 = _8118 | _8115;
    assign _8640 = vdd ? _8119 : gnd;
    assign _7539 = _8640;
    assign _8120 = irq[3:3];
    assign _8121 = _38[3:3];
    assign _8122 = _7536[3:3];
    assign _8123 = _8122 & _8121;
    assign _8124 = _8123 | _8120;
    assign _8639 = vdd ? _8124 : gnd;
    assign _7540 = _8639;
    assign _8125 = irq[4:4];
    assign _8126 = _38[4:4];
    assign _8127 = _7536[4:4];
    assign _8128 = _8127 & _8126;
    assign _8129 = _8128 | _8125;
    assign _8638 = vdd ? _8129 : gnd;
    assign _7541 = _8638;
    assign _8130 = irq[5:5];
    assign _8131 = _38[5:5];
    assign _8132 = _7536[5:5];
    assign _8133 = _8132 & _8131;
    assign _8134 = _8133 | _8130;
    assign _8637 = vdd ? _8134 : gnd;
    assign _7542 = _8637;
    assign _8135 = irq[6:6];
    assign _8136 = _38[6:6];
    assign _8137 = _7536[6:6];
    assign _8138 = _8137 & _8136;
    assign _8139 = _8138 | _8135;
    assign _8636 = vdd ? _8139 : gnd;
    assign _7543 = _8636;
    assign _8140 = irq[7:7];
    assign _8141 = _38[7:7];
    assign _8142 = _7536[7:7];
    assign _8143 = _8142 & _8141;
    assign _8144 = _8143 | _8140;
    assign _8635 = vdd ? _8144 : gnd;
    assign _7544 = _8635;
    assign _8145 = irq[8:8];
    assign _8146 = _38[8:8];
    assign _8147 = _7536[8:8];
    assign _8148 = _8147 & _8146;
    assign _8149 = _8148 | _8145;
    assign _8634 = vdd ? _8149 : gnd;
    assign _7545 = _8634;
    assign _8150 = irq[9:9];
    assign _8151 = _38[9:9];
    assign _8152 = _7536[9:9];
    assign _8153 = _8152 & _8151;
    assign _8154 = _8153 | _8150;
    assign _8633 = vdd ? _8154 : gnd;
    assign _7546 = _8633;
    assign _8155 = irq[10:10];
    assign _8156 = _38[10:10];
    assign _8157 = _7536[10:10];
    assign _8158 = _8157 & _8156;
    assign _8159 = _8158 | _8155;
    assign _8632 = vdd ? _8159 : gnd;
    assign _7547 = _8632;
    assign _8160 = irq[11:11];
    assign _8161 = _38[11:11];
    assign _8162 = _7536[11:11];
    assign _8163 = _8162 & _8161;
    assign _8164 = _8163 | _8160;
    assign _8631 = vdd ? _8164 : gnd;
    assign _7548 = _8631;
    assign _8165 = irq[12:12];
    assign _8166 = _38[12:12];
    assign _8167 = _7536[12:12];
    assign _8168 = _8167 & _8166;
    assign _8169 = _8168 | _8165;
    assign _8630 = vdd ? _8169 : gnd;
    assign _7549 = _8630;
    assign _8170 = irq[13:13];
    assign _8171 = _38[13:13];
    assign _8172 = _7536[13:13];
    assign _8173 = _8172 & _8171;
    assign _8174 = _8173 | _8170;
    assign _8629 = vdd ? _8174 : gnd;
    assign _7550 = _8629;
    assign _8175 = irq[14:14];
    assign _8176 = _38[14:14];
    assign _8177 = _7536[14:14];
    assign _8178 = _8177 & _8176;
    assign _8179 = _8178 | _8175;
    assign _8628 = vdd ? _8179 : gnd;
    assign _7551 = _8628;
    assign _8180 = irq[15:15];
    assign _8181 = _38[15:15];
    assign _8182 = _7536[15:15];
    assign _8183 = _8182 & _8181;
    assign _8184 = _8183 | _8180;
    assign _8627 = vdd ? _8184 : gnd;
    assign _7552 = _8627;
    assign _8185 = irq[16:16];
    assign _8186 = _38[16:16];
    assign _8187 = _7536[16:16];
    assign _8188 = _8187 & _8186;
    assign _8189 = _8188 | _8185;
    assign _8626 = vdd ? _8189 : gnd;
    assign _7553 = _8626;
    assign _8190 = irq[17:17];
    assign _8191 = _38[17:17];
    assign _8192 = _7536[17:17];
    assign _8193 = _8192 & _8191;
    assign _8194 = _8193 | _8190;
    assign _8625 = vdd ? _8194 : gnd;
    assign _7554 = _8625;
    assign _8195 = irq[18:18];
    assign _8196 = _38[18:18];
    assign _8197 = _7536[18:18];
    assign _8198 = _8197 & _8196;
    assign _8199 = _8198 | _8195;
    assign _8624 = vdd ? _8199 : gnd;
    assign _7555 = _8624;
    assign _8200 = irq[19:19];
    assign _8201 = _38[19:19];
    assign _8202 = _7536[19:19];
    assign _8203 = _8202 & _8201;
    assign _8204 = _8203 | _8200;
    assign _8623 = vdd ? _8204 : gnd;
    assign _7556 = _8623;
    assign _8205 = irq[20:20];
    assign _8206 = _38[20:20];
    assign _8207 = _7536[20:20];
    assign _8208 = _8207 & _8206;
    assign _8209 = _8208 | _8205;
    assign _8622 = vdd ? _8209 : gnd;
    assign _7557 = _8622;
    assign _8210 = irq[21:21];
    assign _8211 = _38[21:21];
    assign _8212 = _7536[21:21];
    assign _8213 = _8212 & _8211;
    assign _8214 = _8213 | _8210;
    assign _8621 = vdd ? _8214 : gnd;
    assign _7558 = _8621;
    assign _8215 = irq[22:22];
    assign _8216 = _38[22:22];
    assign _8217 = _7536[22:22];
    assign _8218 = _8217 & _8216;
    assign _8219 = _8218 | _8215;
    assign _8620 = vdd ? _8219 : gnd;
    assign _7559 = _8620;
    assign _8220 = irq[23:23];
    assign _8221 = _38[23:23];
    assign _8222 = _7536[23:23];
    assign _8223 = _8222 & _8221;
    assign _8224 = _8223 | _8220;
    assign _8619 = vdd ? _8224 : gnd;
    assign _7560 = _8619;
    assign _8225 = irq[24:24];
    assign _8226 = _38[24:24];
    assign _8227 = _7536[24:24];
    assign _8228 = _8227 & _8226;
    assign _8229 = _8228 | _8225;
    assign _8618 = vdd ? _8229 : gnd;
    assign _7561 = _8618;
    assign _8230 = irq[25:25];
    assign _8231 = _38[25:25];
    assign _8232 = _7536[25:25];
    assign _8233 = _8232 & _8231;
    assign _8234 = _8233 | _8230;
    assign _8617 = vdd ? _8234 : gnd;
    assign _7562 = _8617;
    assign _8235 = irq[26:26];
    assign _8236 = _38[26:26];
    assign _8237 = _7536[26:26];
    assign _8238 = _8237 & _8236;
    assign _8239 = _8238 | _8235;
    assign _8616 = vdd ? _8239 : gnd;
    assign _7563 = _8616;
    assign _8240 = irq[27:27];
    assign _8241 = _38[27:27];
    assign _8242 = _7536[27:27];
    assign _8243 = _8242 & _8241;
    assign _8244 = _8243 | _8240;
    assign _8615 = vdd ? _8244 : gnd;
    assign _7564 = _8615;
    assign _8245 = irq[28:28];
    assign _8246 = _38[28:28];
    assign _8247 = _7536[28:28];
    assign _8248 = _8247 & _8246;
    assign _8249 = _8248 | _8245;
    assign _8614 = vdd ? _8249 : gnd;
    assign _7565 = _8614;
    assign _8250 = irq[29:29];
    assign _8251 = _38[29:29];
    assign _8252 = _7536[29:29];
    assign _8253 = _8252 & _8251;
    assign _8254 = _8253 | _8250;
    assign _8613 = vdd ? _8254 : gnd;
    assign _7566 = _8613;
    assign _8255 = irq[30:30];
    assign _8256 = _38[30:30];
    assign _8257 = _7536[30:30];
    assign _8258 = _8257 & _8256;
    assign _8259 = _8258 | _8255;
    assign _8612 = vdd ? _8259 : gnd;
    assign _7567 = _8612;
    assign _8260 = irq[31:31];
    assign _8261 = _38[31:31];
    assign _8262 = _7536[31:31];
    assign _8263 = _8262 & _8261;
    assign _8264 = _8263 | _8260;
    assign _8611 = vdd ? _8264 : gnd;
    assign _7568 = _8611;
    assign _7569 = { _7568, _7567, _7566, _7565, _7564, _7563, _7562, _7561, _7560, _7559, _7558, _7557, _7556, _7555, _7554, _7553, _7552, _7551, _7550, _7549, _7548, _7547, _7546, _7545, _7544, _7543, _7542, _7541, _7540, _7539, _7538, _7537 };
    assign _8664 = _6743 == _6740;
    assign _8665 = _8664 ? _8663 : _7569;
    assign _7534 = _8665;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7536 <= _7533;
        else
            _7536 <= _7534;
    end
    assign _9045 = _7536[31:31];
    assign _9046 = _9045 | _9044;
    assign _9047 = _9046 | _9043;
    assign _9048 = _9047 | _9042;
    assign _9049 = _9048 | _9041;
    assign _9050 = _9049 | _9040;
    assign _9051 = _9050 | _9039;
    assign _9052 = _9051 | _9038;
    assign _9053 = _9052 | _9037;
    assign _9054 = _9053 | _9036;
    assign _9055 = _9054 | _9035;
    assign _9056 = _9055 | _9034;
    assign _9057 = _9056 | _9033;
    assign _9058 = _9057 | _9032;
    assign _9059 = _9058 | _9031;
    assign _9060 = _9059 | _9030;
    assign _9061 = _9060 | _9029;
    assign _9062 = _9061 | _9028;
    assign _9063 = _9062 | _9027;
    assign _9064 = _9063 | _9026;
    assign _9065 = _9064 | _9025;
    assign _9066 = _9065 | _9024;
    assign _9067 = _9066 | _9023;
    assign _9068 = _9067 | _9022;
    assign _9069 = _9068 | _9021;
    assign _9070 = _9069 | _9020;
    assign _9071 = _9070 | _9019;
    assign _9072 = _9071 | _9018;
    assign _9073 = _9072 | _9017;
    assign _9074 = _9073 | _9016;
    assign _9075 = _9074 | _9015;
    assign _9076 = _9075 | _9014;
    assign _9077 = _9076 ? _8081 : _7688;
    assign _9078 = _7696 ? _9077 : _8081;
    assign _9079 = _7789 ? _8081 : _9078;
    assign _9080 = _6743 == _6740;
    assign _9081 = _9080 ? _9079 : _8081;
    assign _7470 = _9081;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7472 <= _7469;
        else
            _7472 <= _7470;
    end
    assign _7694 = _6763 | _7472;
    assign _7695 = vdd & _7694;
    assign _7696 = _7695 & _7693;
    assign _8957 = _7696 ? _8956 : _7795;
    assign _8958 = _7789 ? _7795 : _8957;
    assign _8959 = _5634 ? _5637 : _7492;
    assign _8960 = vdd ? _8959 : _7492;
    assign _8961 = vdd ? _8960 : _7492;
    assign _7836 = _5645[46:46];
    assign _7837 = vdd & vdd;
    assign _7838 = _7837 & _7836;
    assign _8962 = _7838 ? _7835 : _7492;
    assign _7873 = _5645[44:44];
    assign _7874 = vdd & _7873;
    assign _8963 = _7874 ? _7872 : _8962;
    assign _8964 = _7880 ? _7875 : _8963;
    assign _8965 = _7886 ? _7881 : _8964;
    assign _8966 = _7890 ? _7887 : _8965;
    assign _8967 = _7894 ? _7492 : _8966;
    assign _8968 = _7910 ? _7895 : _8967;
    assign _8969 = _7925 ? _8961 : _8968;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5821 <= gnd;
        else
            _5821 <= _5769;
    end
    assign _5836 = _5833 ? _5821 : gnd;
    assign _5837 = _5834 ? pcpi_wr : _5836;
    assign _5637 = _5837;
    assign _5811 = _5770 ? vdd : gnd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5721 <= gnd;
        else
            _5721 <= _5719;
    end
    assign _5722 = ~ _5721;
    assign _5688 = _5643[14:12];
    assign _5690 = _5688 == _5689;
    assign _5691 = _5687 & _5690;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5693 <= gnd;
        else
            _5693 <= _5691;
    end
    assign _5712 = _5693 | _5699;
    assign _5713 = _5712 | _5705;
    assign _5714 = _5713 | _5711;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5719 <= gnd;
        else
            _5719 <= _5714;
    end
    assign _5723 = _5719 & _5722;
    assign _5773 = ~ _5723;
    assign _5706 = _5643[14:12];
    assign _5708 = _5706 == _5707;
    assign _5709 = _5687 & _5708;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5711 <= gnd;
        else
            _5711 <= _5709;
    end
    assign _5700 = _5643[14:12];
    assign _5702 = _5700 == _5701;
    assign _5703 = _5687 & _5702;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5705 <= gnd;
        else
            _5705 <= _5703;
    end
    assign _5694 = _5643[14:12];
    assign _5696 = _5694 == _5695;
    assign _5679 = _5643[31:25];
    assign _5681 = _5679 == _5680;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6562 <= _6560;
        else
            if (_5843)
                _6562 <= _5652;
    end
    assign _5643 = _6562;
    assign _5682 = _5643[6:0];
    assign _5684 = _5682 == _5683;
    assign _9295 = _5634 ? _7921 : _7924;
    assign _9296 = vdd ? _9295 : _6767;
    assign _9297 = vdd ? _9296 : _6767;
    assign _9298 = _7925 ? _9297 : _6767;
    assign _9299 = _5634 ? _7936 : _7938;
    assign _9300 = _7940 ? _9299 : _6767;
    assign _9301 = _6743 == _6737;
    assign _9302 = _9301 ? _9300 : _6767;
    assign _9303 = _6743 == _6738;
    assign _9304 = _9303 ? _9298 : _9302;
    assign _6765 = _9304;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6767 <= _6764;
        else
            _6767 <= _6765;
    end
    assign _5665 = _6767;
    assign _5685 = resetn & _5665;
    assign _5686 = _5685 & _5684;
    assign _5687 = _5686 & _5681;
    assign _5697 = _5687 & _5696;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5699 <= gnd;
        else
            _5699 <= _5697;
    end
    assign _5715 = _5699 | _5705;
    assign _5716 = _5715 | _5711;
    assign _5776 = _5716 ? _5775 : _5774;
    assign _5772 = _5763 - _5771;
    assign _5815 = _5766 ? _5776 : _5772;
    assign _5761 = _5815;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5763 <= _5760;
        else
            _5763 <= _5761;
    end
    assign _5770 = _5763[6:6];
    assign _5813 = _5770 ? vdd : _5766;
    assign _5814 = _5766 ? _5773 : _5813;
    assign _5764 = _5814;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5766 <= vdd;
        else
            _5766 <= _5764;
    end
    assign _5812 = _5766 ? gnd : _5811;
    assign _5767 = _5812;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5769 <= gnd;
        else
            _5769 <= _5767;
    end
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5823 <= gnd;
        else
            _5823 <= _5769;
    end
    assign _5833 = vdd & _5823;
    assign _5834 = gnd & pcpi_ready;
    assign _5835 = _5834 | _5833;
    assign _5634 = _5835;
    assign _8970 = _5634 ? _5637 : _7492;
    assign _7939 = _5645[47:47];
    assign _7940 = vdd & _7939;
    assign _8971 = _7940 ? _8970 : _7492;
    assign _8972 = _7948 ? _7422 : _7943;
    assign _8973 = _6743 == _6733;
    assign _8974 = _8973 ? _8073 : _7492;
    assign _8975 = _6743 == _6735;
    assign _8976 = _8975 ? _8006 : _8974;
    assign _8977 = _6743 == _6736;
    assign _8978 = _8977 ? _8972 : _8976;
    assign _8979 = _6743 == _6737;
    assign _8980 = _8979 ? _8971 : _8978;
    assign _8981 = _6743 == _6738;
    assign _8982 = _8981 ? _8969 : _8980;
    assign _8983 = _6743 == _6740;
    assign _8984 = _8983 ? _8958 : _8982;
    assign _7490 = _8984;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7492 <= _7489;
        else
            _7492 <= _7490;
    end
    assign _8667 = _7492 ? _7532 : _8666;
    assign _8668 = _7484 ? _7532 : _8667;
    assign _8669 = _7880 ? _7877 : _7532;
    assign _8670 = _7886 ? _7532 : _8669;
    assign _8671 = _7890 ? _7532 : _8670;
    assign _8672 = _7894 ? _7532 : _8671;
    assign _8673 = _7910 ? _7532 : _8672;
    assign _8674 = _7925 ? _7532 : _8673;
    assign _8675 = _6743 == _6738;
    assign _8676 = _8675 ? _8674 : _7532;
    assign _8677 = _6743 == _6740;
    assign _8678 = _8677 ? _8668 : _8676;
    assign _7530 = _8678;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7532 <= _7529;
        else
            _7532 <= _7530;
    end
    assign _7785 = ~ _7532;
    assign _7786 = _6763 & _7785;
    assign _7787 = _7786 & _7784;
    assign _7788 = _7787 | _7719;
    assign _7789 = vdd & _7788;
    assign _8993 = _7789 ? _7793 : _8992;
    assign _7879 = _5645[43:43];
    assign _7880 = vdd & _7879;
    assign _8994 = _7880 ? _7876 : _7484;
    assign _7884 = _5645[42:42];
    assign _7885 = vdd & vdd;
    assign _7886 = _7885 & _7884;
    assign _8995 = _7886 ? _7484 : _8994;
    assign _7888 = _5645[41:41];
    assign _7889 = vdd & vdd;
    assign _7890 = _7889 & _7888;
    assign _8996 = _7890 ? _7484 : _8995;
    assign _7894 = _5644[0:0];
    assign _8997 = _7894 ? _7484 : _8996;
    assign _7910 = _5644[14:14];
    assign _8998 = _7910 ? _7484 : _8997;
    assign _7925 = _5645[47:47];
    assign _8999 = _7925 ? _7484 : _8998;
    assign _7944 = _5645[3:3];
    assign _9000 = _7948 ? _7422 : _7944;
    assign _9001 = _6743 == _6736;
    assign _9002 = _9001 ? _9000 : _7484;
    assign _9003 = _6743 == _6738;
    assign _9004 = _9003 ? _8999 : _9002;
    assign _9005 = _6743 == _6740;
    assign _9006 = _9005 ? _8993 : _9004;
    assign _7482 = _9006;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7484 <= _7481;
        else
            _7484 <= _7482;
    end
    assign _9110 = _7484 ? _9103 : _9109;
    assign _9111 = _6743 == _6740;
    assign _9112 = _9111 ? _9110 : _6808;
    assign _6809 = _9112;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7205 <= _7203;
        else
            if (_7202)
                _7205 <= _6809;
    end
    always @* begin
        case (_5640)
        0: _7381 <= _7205;
        1: _7381 <= _7210;
        2: _7381 <= _7215;
        3: _7381 <= _7220;
        4: _7381 <= _7225;
        5: _7381 <= _7230;
        6: _7381 <= _7235;
        7: _7381 <= _7240;
        8: _7381 <= _7245;
        9: _7381 <= _7250;
        10: _7381 <= _7255;
        11: _7381 <= _7260;
        12: _7381 <= _7265;
        13: _7381 <= _7270;
        14: _7381 <= _7275;
        15: _7381 <= _7280;
        16: _7381 <= _7285;
        17: _7381 <= _7290;
        18: _7381 <= _7295;
        19: _7381 <= _7300;
        20: _7381 <= _7305;
        21: _7381 <= _7310;
        22: _7381 <= _7315;
        23: _7381 <= _7320;
        24: _7381 <= _7325;
        25: _7381 <= _7330;
        26: _7381 <= _7335;
        27: _7381 <= _7340;
        28: _7381 <= _7345;
        29: _7381 <= _7350;
        30: _7381 <= _7355;
        31: _7381 <= _7360;
        32: _7381 <= _7365;
        33: _7381 <= _7370;
        34: _7381 <= _7375;
        default: _7381 <= _7380;
        endcase
    end
    assign _6547 = _5653[24:20];
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6550 <= _6548;
        else
            if (_5841)
                _6550 <= _6547;
    end
    assign _6551 = { gnd, _6550 };
    assign _5640 = _6551;
    assign _7823 = _5640 == _7822;
    assign _7824 = ~ _7823;
    assign _7825 = _7824 ? _7381 : _7821;
    assign _7941 = _7825[4:0];
    assign _7975 = _7524 - _7974;
    assign _7951 = _7524 - _7950;
    assign _8002 = _7524 < _8001;
    assign _8003 = ~ _8002;
    assign _8696 = _8003 ? _7975 : _7951;
    assign _8697 = _8005 ? _8266 : _8696;
    assign _8698 = _6743 == _6735;
    assign _8699 = _8698 ? _8697 : _8266;
    assign _8700 = _6743 == _6737;
    assign _8701 = _8700 ? _7941 : _8699;
    assign _8702 = _6743 == _6738;
    assign _8703 = _8702 ? _8695 : _8701;
    assign _7522 = _8703;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7524 <= _7521;
        else
            _7524 <= _7522;
    end
    assign _8005 = _7524 == _8004;
    assign _9138 = _8005 ? _6799 : _9137;
    assign _8012 = _6799 + _5639;
    assign _9139 = _8023 ? _8012 : _6799;
    assign _9140 = _8025 ? _9139 : _6799;
    assign _9317 = _8010 ? _8007 : _8082;
    assign _9318 = _8025 ? _9317 : _8082;
    assign _9319 = _8050 ? _8026 : _8082;
    assign _9320 = _8072 ? _9319 : _8082;
    assign _9321 = _6743 == _6733;
    assign _9322 = _9321 ? _9320 : _8082;
    assign _9323 = _6743 == _6734;
    assign _9324 = _9323 ? _9318 : _9322;
    assign _6753 = _9324;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6755 <= _6752;
        else
            _6755 <= _6753;
    end
    assign _5662 = _6755;
    assign _5842 = ~ _5662;
    assign _5843 = _5664 & _5842;
    assign _5841 = _5670 & _5659;
    assign _6485 = _6480[0:0];
    assign _6482 = _6480[19:10];
    assign _6483 = _6480[9:9];
    assign _6484 = _6480[8:1];
    assign _6475 = { _6474, _6473 };
    assign _6471 = _5653[31:12];
    assign _6472 = { _6471, gnd };
    assign _6473 = _6472[20:20];
    assign _6474 = { _6473, _6473 };
    assign _6476 = { _6474, _6474 };
    assign _6477 = { _6476, _6476 };
    assign _6478 = { _6477, _6475 };
    assign _6480 = { _6478, _6472 };
    assign _6481 = _6480[31:20];
    assign _6486 = { _6481, _6484, _6483, _6482, _6485 };
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6489 <= _6487;
        else
            if (_5841)
                _6489 <= _6486;
    end
    assign _6533 = _5652[31:12];
    assign _6534 = { _6533, _6532 };
    assign _6518 = _5652[31:20];
    assign _6519 = _6518[11:11];
    assign _6520 = { _6519, _6519 };
    assign _6521 = { _6520, _6520 };
    assign _6522 = { _6521, _6521 };
    assign _6523 = { _6522, _6522 };
    assign _6524 = { _6523, _6521 };
    assign _6526 = { _6524, _6518 };
    assign _6510 = { _6509, _6508 };
    assign _6506 = _5652[11:8];
    assign _6505 = _5652[30:25];
    assign _6504 = _5652[7:7];
    assign _6503 = _5652[31:31];
    assign _6507 = { _6503, _6504, _6505, _6506, gnd };
    assign _6508 = _6507[12:12];
    assign _6509 = { _6508, _6508 };
    assign _6511 = { _6509, _6509 };
    assign _6512 = { _6511, _6511 };
    assign _6513 = { _6512, _6512 };
    assign _6514 = { _6513, _6510 };
    assign _6516 = { _6514, _6507 };
    assign _6492 = _5652[11:7];
    assign _6491 = _5652[31:25];
    assign _6493 = { _6491, _6492 };
    assign _6494 = _6493[11:11];
    assign _6495 = { _6494, _6494 };
    assign _6496 = { _6495, _6495 };
    assign _6497 = { _6496, _6496 };
    assign _6498 = { _6497, _6497 };
    assign _6499 = { _6498, _6496 };
    assign _6501 = { _6499, _6493 };
    assign _6502 = _6446[4:4];
    assign _6539 = _6502 ? _6501 : _6490;
    assign _6517 = _6446[9:9];
    assign _6540 = _6517 ? _6516 : _6539;
    assign _6528 = _6446[11:11];
    assign _6527 = _6446[1:1];
    assign _6529 = _6527 | _6528;
    assign _6530 = _6308[3:3];
    assign _6531 = _6530 | _6529;
    assign _6541 = _6531 ? _6526 : _6540;
    assign _6536 = _6308[1:1];
    assign _6535 = _6308[0:0];
    assign _6537 = _6535 | _6536;
    assign _6542 = _6537 ? _6534 : _6541;
    assign _6538 = _6308[2:2];
    assign _6543 = _6538 ? _6489 : _6542;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6546 <= _6544;
        else
            if (_5843)
                _6546 <= _6543;
    end
    assign _5639 = _6546;
    assign _8052 = _6799 + _5639;
    assign _9141 = _8070 ? _8052 : _6799;
    assign _9142 = _8072 ? _9141 : _6799;
    assign _9143 = _6743 == _6733;
    assign _9144 = _9143 ? _9142 : _6799;
    assign _9145 = _6743 == _6734;
    assign _9146 = _9145 ? _9140 : _9144;
    assign _9147 = _6743 == _6735;
    assign _9148 = _9147 ? _9138 : _9146;
    assign _9149 = _6743 == _6738;
    assign _9150 = _9149 ? _9136 : _9148;
    assign _6797 = _9150;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6799 <= _6796;
        else
            _6799 <= _6797;
    end
    assign _7383 = _6799 < _6795;
    assign _7394 = _5644[7:7];
    assign _7414 = _7394 ? _7393 : _7383;
    assign _7397 = _5645[9:9];
    assign _7408 = _5645[7:7];
    assign _7417 = _7408 | _7397;
    assign _7411 = _5645[5:5];
    assign _5645 = _6308;
    assign _7413 = _5645[4:4];
    assign _7419 = _7413 | _7411;
    assign _7421 = _7419 | _7417;
    assign _7422 = _7421 ? _7420 : _7414;
    assign _9305 = _7422 ? _7946 : _8083;
    assign _9306 = _7948 ? _9305 : _8083;
    assign _8009 = ~ _6771;
    assign _8010 = _8009 & _5659;
    assign _9307 = _8010 ? _8008 : _8083;
    assign _9308 = _8025 ? _9307 : _8083;
    assign _8049 = ~ _6771;
    assign _8050 = _8049 & _5659;
    assign _9309 = _8050 ? _8027 : _8083;
    assign _9310 = _8072 ? _9309 : _8083;
    assign _8083 = _6787 & _5659;
    assign _9311 = _6743 == _6733;
    assign _9312 = _9311 ? _9310 : _8083;
    assign _9313 = _6743 == _6734;
    assign _9314 = _9313 ? _9308 : _9312;
    assign _9315 = _6743 == _6736;
    assign _9316 = _9315 ? _9306 : _9314;
    assign _6761 = _9316;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6763 <= _6760;
        else
            _6763 <= _6761;
    end
    assign _5664 = _6763;
    assign _5846 = _5664 & _5845;
    assign _5652 = _6602;
    assign _6235 = _5652[14:12];
    assign _6237 = _6235 == _6236;
    assign _5867 = _5653[6:0];
    assign _5869 = _5867 == _5868;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_beq_bne_blt_bge_bltu_bgeu <= gnd;
        else
            if (_5844)
                is_beq_bne_blt_bge_bltu_bgeu <= _5869;
    end
    assign _6238 = is_beq_bne_blt_bge_bltu_bgeu & _6237;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_beq <= gnd;
        else
            if (_5846)
                instr_beq <= _6238;
    end
    assign _6241 = _5653[31:25];
    assign _6243 = _6241 == _6242;
    assign _6244 = _5653[6:0];
    assign _6246 = _6244 == _6245;
    assign _6247 = _6246 & _6243;
    assign _6248 = _6247 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_waitirq <= gnd;
        else
            if (_5844)
                instr_waitirq <= _6248;
    end
    assign _6251 = _5653[31:25];
    assign _6253 = _6251 == _6252;
    assign _6254 = _5653[6:0];
    assign _6256 = _6254 == _6255;
    assign _6257 = _6256 & _6253;
    assign _6258 = _6257 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_retirq <= gnd;
        else
            if (_5844)
                instr_retirq <= _6258;
    end
    assign _5862 = _5653[6:0];
    assign _5864 = _5862 == _5863;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_jalr <= gnd;
        else
            if (_5844)
                instr_jalr <= _5864;
    end
    assign _5857 = _5653[6:0];
    assign _5859 = _5857 == _5858;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_jal <= gnd;
        else
            if (_5844)
                instr_jal <= _5859;
    end
    assign _5852 = _5653[6:0];
    assign _5854 = _5852 == _5853;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_auipc <= gnd;
        else
            if (_5844)
                instr_auipc <= _5854;
    end
    assign _5844 = _5670 & _5659;
    assign _6599 = _6577 & mem_ready;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6602 <= _6600;
        else
            if (_6599)
                _6602 <= _6598;
    end
    assign _9276 = _5659 ? _8078 : _6779;
    assign _8070 = ~ _6779;
    assign _8283 = _8070 ? _8051 : gnd;
    assign _8284 = _8072 ? _8283 : gnd;
    assign _8285 = _6743 == _6733;
    assign _8286 = _8285 ? _8284 : gnd;
    assign _7668 = _8286;
    assign _9277 = _7668 ? _8075 : _9276;
    assign _6777 = _9277;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6779 <= _6776;
        else
            _6779 <= _6777;
    end
    assign _5668 = _6779;
    assign _5666 = _6771;
    assign _6695 = _5666 | _5670;
    assign _6696 = _6695 | _5668;
    assign _6708 = _6696 ? vdd : _6577;
    assign _9274 = _5659 ? _8077 : _6783;
    assign _8023 = ~ _6783;
    assign _8287 = _8023 ? _8011 : gnd;
    assign _8024 = ~ _6771;
    assign _8025 = _8024 | _5659;
    assign _8288 = _8025 ? _8287 : gnd;
    assign _8289 = _6743 == _6734;
    assign _8290 = _8289 ? _8288 : gnd;
    assign _7667 = _8290;
    assign _9275 = _7667 ? _8074 : _9274;
    assign _6781 = _9275;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6783 <= _6780;
        else
            _6783 <= _6781;
    end
    assign _5669 = _6783;
    assign _6709 = _5669 ? vdd : _6708;
    assign _6710 = mem_ready ? gnd : _6577;
    assign _6711 = mem_ready ? gnd : _6577;
    assign _6712 = _6570 == _6565;
    assign _6713 = _6712 ? _6711 : _6577;
    assign _6714 = _6570 == _6566;
    assign _6715 = _6714 ? _6710 : _6713;
    assign _6716 = _6570 == _6567;
    assign _6717 = _6716 ? _6709 : _6715;
    assign _6575 = _6717;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6577 <= gnd;
        else
            _6577 <= _6575;
    end
    assign _6603 = _6577 & mem_ready;
    assign _6604 = _6603 | gnd;
    assign _6605 = _6604 ? mem_rdata : _6602;
    assign _6598 = _6605;
    assign _5653 = _6598;
    assign _5847 = _5653[6:0];
    assign _5849 = _5847 == _5848;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lui <= gnd;
        else
            if (_5844)
                instr_lui <= _5849;
    end
    assign _6261 = instr_lui | instr_auipc;
    assign _6262 = _6261 | instr_jal;
    assign _6263 = _6262 | instr_jalr;
    assign _6264 = _6263 | instr_retirq;
    assign _6265 = _6264 | instr_waitirq;
    assign _6266 = _6265 | instr_beq;
    assign _6267 = _6266 | instr_bne;
    assign _6268 = _6267 | instr_blt;
    assign _6269 = _6268 | instr_bge;
    assign _6270 = _6269 | instr_bltu;
    assign _6271 = _6270 | instr_bgeu;
    assign _6272 = _6271 | instr_lb;
    assign _6273 = _6272 | instr_lh;
    assign _6274 = _6273 | instr_lw;
    assign _6275 = _6274 | instr_lbu;
    assign _6276 = _6275 | instr_lhu;
    assign _6277 = _6276 | instr_sb;
    assign _6278 = _6277 | instr_sh;
    assign _6279 = _6278 | instr_sw;
    assign _6280 = _6279 | instr_addi;
    assign _6281 = _6280 | instr_slti;
    assign _6282 = _6281 | instr_sltiu;
    assign _6283 = _6282 | instr_xori;
    assign _6284 = _6283 | instr_ori;
    assign _6285 = _6284 | instr_andi;
    assign _6286 = _6285 | instr_slli;
    assign _6287 = _6286 | instr_srli;
    assign _6288 = _6287 | instr_srai;
    assign _6289 = _6288 | instr_add;
    assign _6290 = _6289 | instr_sub;
    assign _6291 = _6290 | instr_sll;
    assign _6292 = _6291 | instr_slt;
    assign _6293 = _6292 | instr_sltu;
    assign _6294 = _6293 | instr_xor;
    assign _6295 = _6294 | instr_srl;
    assign _6296 = _6295 | instr_sra;
    assign _6297 = _6296 | instr_or;
    assign _6298 = _6297 | instr_and;
    assign _6299 = _6298 | instr_rdcycle;
    assign _6300 = _6299 | instr_rdcycleh;
    assign _6301 = _6300 | instr_rdinstr;
    assign _6302 = _6301 | instr_rdinstrh;
    assign _6303 = _6302 | instr_getq;
    assign _6304 = _6303 | instr_setq;
    assign _6305 = _6304 | instr_maskirq;
    assign _6306 = _6305 | instr_timer;
    assign instr_trap = ~ _6306;
    assign _6308 = { instr_trap, instr_timer, instr_waitirq, instr_maskirq, instr_retirq, instr_setq, instr_getq, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle, instr_and, instr_or, instr_sra, instr_srl, instr_xor, instr_sltu, instr_slt, instr_sll, instr_sub, instr_add, instr_srai, instr_srli, instr_slli, instr_andi, instr_ori, instr_xori, instr_sltiu, instr_slti, instr_addi, instr_sw, instr_sh, instr_sb, instr_lhu, instr_lbu, instr_lw, instr_lh, instr_lb, instr_bgeu, instr_bltu, instr_bge, instr_blt, instr_bne, instr_beq, instr_jalr, instr_jal, instr_auipc, instr_lui };
    assign _6309 = _6308[37:37];
    assign _6313 = _6309 | _6310;
    assign _6314 = _6313 | _6311;
    assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = _6314 | _6312;
    assign _6446 = { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_compare, is_alu_reg_reg, is_alu_reg_imm, is_lbu_lhu_lw, is_beq_bne_blt_bge_bltu_bgeu, is_sltiu_bltu_sltu, is_slti_blt_slt, is_lui_auipc_jal_jalr_addi_add, is_sll_srl_sra, is_sb_sh_sw, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lb_lh_lw_lbu_lhu, is_lui_auipc_jal };
    assign _5644 = _6446;
    assign _7948 = _5644[9:9];
    assign _8280 = _7948 ? _8279 : gnd;
    assign _8281 = _6743 == _6736;
    assign _8282 = _8281 ? _8280 : gnd;
    assign _7669 = _8282;
    assign _9273 = _7669 ? _8076 : _9272;
    assign _6785 = _9273;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6787 <= _6784;
        else
            _6787 <= _6785;
    end
    assign _5670 = _6787;
    assign _6723 = _5670 ? _6567 : _6570;
    assign _6724 = _6570 == _6564;
    assign _6725 = _6724 ? _6723 : _6570;
    assign _6726 = _6570 == _6565;
    assign _6727 = _6726 ? _6722 : _6725;
    assign _6728 = _6570 == _6566;
    assign _6729 = _6728 ? _6721 : _6727;
    assign _6730 = _6570 == _6567;
    assign _6731 = _6730 ? _6719 : _6729;
    assign _6568 = _6731;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6570 <= _6563;
        else
            _6570 <= _6568;
    end
    assign _6573 = _6567 == _6570;
    assign _6574 = ~ _6573;
    assign _6584 = mem_ready & _6574;
    assign _6585 = _6584 & _6583;
    assign _6586 = _6585 | _6581;
    assign _5659 = _6586;
    assign _9294 = _5659 ? _8080 : _9293;
    assign _6769 = _9294;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6771 <= _6768;
        else
            _6771 <= _6769;
    end
    assign _8071 = ~ _6771;
    assign _8072 = _8071 | _5659;
    assign _9375 = _8072 ? _9374 : _6743;
    assign _9376 = _6743 == _6733;
    assign _9377 = _9376 ? _9375 : _6743;
    assign _9378 = _6743 == _6734;
    assign _9379 = _9378 ? _9373 : _9377;
    assign _9380 = _6743 == _6735;
    assign _9381 = _9380 ? _9371 : _9379;
    assign _9382 = _6743 == _6736;
    assign _9383 = _9382 ? _9370 : _9381;
    assign _9384 = _6743 == _6737;
    assign _9385 = _9384 ? _9368 : _9383;
    assign _9386 = _6743 == _6738;
    assign _9387 = _9386 ? _9362 : _9385;
    assign _9388 = _6743 == _6740;
    assign _9389 = _9388 ? _9342 : _9387;
    assign _6741 = _9389;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6743 <= _6732;
        else
            _6743 <= _6741;
    end
    assign _9169 = _6743 == _6739;
    assign _9170 = _9169 ? vdd : _8267;
    assign _6789 = _9170;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6791 <= _6788;
        else
            _6791 <= _6789;
    end
    assign _5671 = _6791;

    /* aliases */

    /* output assignments */
    assign trap = _5671;
    assign mem_valid = _5658;
    assign mem_instr = _5657;
    assign mem_addr = _5656;
    assign mem_wdata = _5655;
    assign mem_wstrb = _5654;
    assign mem_la_read = _5650;
    assign mem_la_write = _5649;
    assign mem_la_addr = _5648;
    assign mem_la_wdata = _5647;
    assign mem_la_wstrb = _5646;
    assign pcpi_valid = _5665;
    assign pcpi_insn = _5643;
    assign pcpi_rs1 = _5673;
    assign pcpi_rs2 = _5672;
    assign eoi = _5661;

endmodule
