module opicorv32_rf (
    ra2,
    wa,
    wr,
    resetn,
    clk,
    d,
    ra1,
    q1,
    q2
);

    input [5:0] ra2;
    input [5:0] wa;
    input wr;
    input resetn;
    input clk;
    input [31:0] d;
    input [5:0] ra1;
    output [31:0] q1;
    output [31:0] q2;

    /* signal declarations */
    reg [31:0] _2342;
    wire _2337;
    wire _2338;
    wire [31:0] _2340 = 32'b00000000000000000000000000000000;
    wire [31:0] _2339 = 32'b00000000000000000000000000000000;
    reg [31:0] _2341;
    wire _2332;
    wire _2333;
    wire [31:0] _2335 = 32'b00000000000000000000000000000000;
    wire [31:0] _2334 = 32'b00000000000000000000000000000000;
    reg [31:0] _2336;
    wire _2327;
    wire _2328;
    wire [31:0] _2330 = 32'b00000000000000000000000000000000;
    wire [31:0] _2329 = 32'b00000000000000000000000000000000;
    reg [31:0] _2331;
    wire _2322;
    wire _2323;
    wire [31:0] _2325 = 32'b00000000000000000000000000000000;
    wire [31:0] _2324 = 32'b00000000000000000000000000000000;
    reg [31:0] _2326;
    wire _2317;
    wire _2318;
    wire [31:0] _2320 = 32'b00000000000000000000000000000000;
    wire [31:0] _2319 = 32'b00000000000000000000000000000000;
    reg [31:0] _2321;
    wire _2312;
    wire _2313;
    wire [31:0] _2315 = 32'b00000000000000000000000000000000;
    wire [31:0] _2314 = 32'b00000000000000000000000000000000;
    reg [31:0] _2316;
    wire _2307;
    wire _2308;
    wire [31:0] _2310 = 32'b00000000000000000000000000000000;
    wire [31:0] _2309 = 32'b00000000000000000000000000000000;
    reg [31:0] _2311;
    wire _2302;
    wire _2303;
    wire [31:0] _2305 = 32'b00000000000000000000000000000000;
    wire [31:0] _2304 = 32'b00000000000000000000000000000000;
    reg [31:0] _2306;
    wire _2297;
    wire _2298;
    wire [31:0] _2300 = 32'b00000000000000000000000000000000;
    wire [31:0] _2299 = 32'b00000000000000000000000000000000;
    reg [31:0] _2301;
    wire _2292;
    wire _2293;
    wire [31:0] _2295 = 32'b00000000000000000000000000000000;
    wire [31:0] _2294 = 32'b00000000000000000000000000000000;
    reg [31:0] _2296;
    wire _2287;
    wire _2288;
    wire [31:0] _2290 = 32'b00000000000000000000000000000000;
    wire [31:0] _2289 = 32'b00000000000000000000000000000000;
    reg [31:0] _2291;
    wire _2282;
    wire _2283;
    wire [31:0] _2285 = 32'b00000000000000000000000000000000;
    wire [31:0] _2284 = 32'b00000000000000000000000000000000;
    reg [31:0] _2286;
    wire _2277;
    wire _2278;
    wire [31:0] _2280 = 32'b00000000000000000000000000000000;
    wire [31:0] _2279 = 32'b00000000000000000000000000000000;
    reg [31:0] _2281;
    wire _2272;
    wire _2273;
    wire [31:0] _2275 = 32'b00000000000000000000000000000000;
    wire [31:0] _2274 = 32'b00000000000000000000000000000000;
    reg [31:0] _2276;
    wire _2267;
    wire _2268;
    wire [31:0] _2270 = 32'b00000000000000000000000000000000;
    wire [31:0] _2269 = 32'b00000000000000000000000000000000;
    reg [31:0] _2271;
    wire _2262;
    wire _2263;
    wire [31:0] _2265 = 32'b00000000000000000000000000000000;
    wire [31:0] _2264 = 32'b00000000000000000000000000000000;
    reg [31:0] _2266;
    wire _2257;
    wire _2258;
    wire [31:0] _2260 = 32'b00000000000000000000000000000000;
    wire [31:0] _2259 = 32'b00000000000000000000000000000000;
    reg [31:0] _2261;
    wire _2252;
    wire _2253;
    wire [31:0] _2255 = 32'b00000000000000000000000000000000;
    wire [31:0] _2254 = 32'b00000000000000000000000000000000;
    reg [31:0] _2256;
    wire _2247;
    wire _2248;
    wire [31:0] _2250 = 32'b00000000000000000000000000000000;
    wire [31:0] _2249 = 32'b00000000000000000000000000000000;
    reg [31:0] _2251;
    wire _2242;
    wire _2243;
    wire [31:0] _2245 = 32'b00000000000000000000000000000000;
    wire [31:0] _2244 = 32'b00000000000000000000000000000000;
    reg [31:0] _2246;
    wire _2237;
    wire _2238;
    wire [31:0] _2240 = 32'b00000000000000000000000000000000;
    wire [31:0] _2239 = 32'b00000000000000000000000000000000;
    reg [31:0] _2241;
    wire _2232;
    wire _2233;
    wire [31:0] _2235 = 32'b00000000000000000000000000000000;
    wire [31:0] _2234 = 32'b00000000000000000000000000000000;
    reg [31:0] _2236;
    wire _2227;
    wire _2228;
    wire [31:0] _2230 = 32'b00000000000000000000000000000000;
    wire [31:0] _2229 = 32'b00000000000000000000000000000000;
    reg [31:0] _2231;
    wire _2222;
    wire _2223;
    wire [31:0] _2225 = 32'b00000000000000000000000000000000;
    wire [31:0] _2224 = 32'b00000000000000000000000000000000;
    reg [31:0] _2226;
    wire _2217;
    wire _2218;
    wire [31:0] _2220 = 32'b00000000000000000000000000000000;
    wire [31:0] _2219 = 32'b00000000000000000000000000000000;
    reg [31:0] _2221;
    wire _2212;
    wire _2213;
    wire [31:0] _2215 = 32'b00000000000000000000000000000000;
    wire [31:0] _2214 = 32'b00000000000000000000000000000000;
    reg [31:0] _2216;
    wire _2207;
    wire _2208;
    wire [31:0] _2210 = 32'b00000000000000000000000000000000;
    wire [31:0] _2209 = 32'b00000000000000000000000000000000;
    reg [31:0] _2211;
    wire _2202;
    wire _2203;
    wire [31:0] _2205 = 32'b00000000000000000000000000000000;
    wire [31:0] _2204 = 32'b00000000000000000000000000000000;
    reg [31:0] _2206;
    wire _2197;
    wire _2198;
    wire [31:0] _2200 = 32'b00000000000000000000000000000000;
    wire [31:0] _2199 = 32'b00000000000000000000000000000000;
    reg [31:0] _2201;
    wire _2192;
    wire _2193;
    wire [31:0] _2195 = 32'b00000000000000000000000000000000;
    wire [31:0] _2194 = 32'b00000000000000000000000000000000;
    reg [31:0] _2196;
    wire _2187;
    wire _2188;
    wire [31:0] _2190 = 32'b00000000000000000000000000000000;
    wire [31:0] _2189 = 32'b00000000000000000000000000000000;
    reg [31:0] _2191;
    wire _2182;
    wire _2183;
    wire [31:0] _2185 = 32'b00000000000000000000000000000000;
    wire [31:0] _2184 = 32'b00000000000000000000000000000000;
    reg [31:0] _2186;
    wire _2177;
    wire _2178;
    wire [31:0] _2180 = 32'b00000000000000000000000000000000;
    wire [31:0] _2179 = 32'b00000000000000000000000000000000;
    reg [31:0] _2181;
    wire _2172;
    wire _2173;
    wire [31:0] _2175 = 32'b00000000000000000000000000000000;
    wire [31:0] _2174 = 32'b00000000000000000000000000000000;
    reg [31:0] _2176;
    wire _2167;
    wire _2168;
    wire [31:0] _2170 = 32'b00000000000000000000000000000000;
    wire [31:0] _2169 = 32'b00000000000000000000000000000000;
    reg [31:0] _2171;
    wire _1778;
    wire _1781;
    wire _1789;
    wire _1809;
    wire _1857;
    wire _1969;
    wire _1779;
    wire _1780;
    wire _1788;
    wire _1808;
    wire _1856;
    wire _1968;
    wire _1782;
    wire _1784;
    wire _1787;
    wire _1807;
    wire _1855;
    wire _1967;
    wire _1783;
    wire _1785;
    wire _1786;
    wire _1806;
    wire _1854;
    wire _1966;
    wire _1790;
    wire _1793;
    wire _1800;
    wire _1805;
    wire _1853;
    wire _1965;
    wire _1791;
    wire _1792;
    wire _1799;
    wire _1804;
    wire _1852;
    wire _1964;
    wire _1794;
    wire _1796;
    wire _1798;
    wire _1803;
    wire _1851;
    wire _1963;
    wire _1795;
    wire _1797;
    wire _1801;
    wire _1802;
    wire _1850;
    wire _1962;
    wire _1810;
    wire _1813;
    wire _1821;
    wire _1840;
    wire _1849;
    wire _1961;
    wire _1811;
    wire _1812;
    wire _1820;
    wire _1839;
    wire _1848;
    wire _1960;
    wire _1814;
    wire _1816;
    wire _1819;
    wire _1838;
    wire _1847;
    wire _1959;
    wire _1815;
    wire _1817;
    wire _1818;
    wire _1837;
    wire _1846;
    wire _1958;
    wire _1822;
    wire _1825;
    wire _1832;
    wire _1836;
    wire _1845;
    wire _1957;
    wire _1823;
    wire _1824;
    wire _1831;
    wire _1835;
    wire _1844;
    wire _1956;
    wire _1826;
    wire _1828;
    wire _1830;
    wire _1834;
    wire _1843;
    wire _1955;
    wire _1827;
    wire _1829;
    wire _1833;
    wire _1841;
    wire _1842;
    wire _1954;
    wire _1858;
    wire _1861;
    wire _1869;
    wire _1889;
    wire _1936;
    wire _1953;
    wire _1859;
    wire _1860;
    wire _1868;
    wire _1888;
    wire _1935;
    wire _1952;
    wire _1862;
    wire _1864;
    wire _1867;
    wire _1887;
    wire _1934;
    wire _1951;
    wire _1863;
    wire _1865;
    wire _1866;
    wire _1886;
    wire _1933;
    wire _1950;
    wire _1870;
    wire _1873;
    wire _1880;
    wire _1885;
    wire _1932;
    wire _1949;
    wire _1871;
    wire _1872;
    wire _1879;
    wire _1884;
    wire _1931;
    wire _1948;
    wire _1874;
    wire _1876;
    wire _1878;
    wire _1883;
    wire _1930;
    wire _1947;
    wire _1875;
    wire _1877;
    wire _1881;
    wire _1882;
    wire _1929;
    wire _1946;
    wire _1890;
    wire _1893;
    wire _1901;
    wire _1920;
    wire _1928;
    wire _1945;
    wire _1891;
    wire _1892;
    wire _1900;
    wire _1919;
    wire _1927;
    wire _1944;
    wire _1894;
    wire _1896;
    wire _1899;
    wire _1918;
    wire _1926;
    wire _1943;
    wire _1895;
    wire _1897;
    wire _1898;
    wire _1917;
    wire _1925;
    wire _1942;
    wire _1902;
    wire _1905;
    wire _1912;
    wire _1916;
    wire _1924;
    wire _1941;
    wire _1903;
    wire _1904;
    wire _1911;
    wire _1915;
    wire _1923;
    wire _1940;
    wire _1906;
    wire _1908;
    wire _1910;
    wire _1914;
    wire _1922;
    wire _1939;
    wire _1907;
    wire _1909;
    wire _1913;
    wire _1921;
    wire _1937;
    wire _1938;
    wire _1970;
    wire _1973;
    wire _1981;
    wire _2001;
    wire _2049;
    wire _2160;
    wire _1971;
    wire _1972;
    wire _1980;
    wire _2000;
    wire _2048;
    wire _2159;
    wire _1974;
    wire _1976;
    wire _1979;
    wire _1999;
    wire _2047;
    wire _2158;
    wire _1975;
    wire _1977;
    wire _1978;
    wire _1998;
    wire _2046;
    wire _2157;
    wire _1982;
    wire _1985;
    wire _1992;
    wire _1997;
    wire _2045;
    wire _2156;
    wire _1983;
    wire _1984;
    wire _1991;
    wire _1996;
    wire _2044;
    wire _2155;
    wire _1986;
    wire _1988;
    wire _1990;
    wire _1995;
    wire _2043;
    wire _2154;
    wire _1987;
    wire _1989;
    wire _1993;
    wire _1994;
    wire _2042;
    wire _2153;
    wire _2002;
    wire _2005;
    wire _2013;
    wire _2032;
    wire _2041;
    wire _2152;
    wire _2003;
    wire _2004;
    wire _2012;
    wire _2031;
    wire _2040;
    wire _2151;
    wire _2006;
    wire _2008;
    wire _2011;
    wire _2030;
    wire _2039;
    wire _2150;
    wire _2007;
    wire _2009;
    wire _2010;
    wire _2029;
    wire _2038;
    wire _2149;
    wire _2014;
    wire _2017;
    wire _2024;
    wire _2028;
    wire _2037;
    wire _2148;
    wire _2015;
    wire _2016;
    wire _2023;
    wire _2027;
    wire _2036;
    wire _2147;
    wire _2018;
    wire _2020;
    wire _2022;
    wire _2026;
    wire _2035;
    wire _2146;
    wire _2019;
    wire _2021;
    wire _2025;
    wire _2033;
    wire _2034;
    wire _2145;
    wire _2050;
    wire _2053;
    wire _2061;
    wire _2081;
    wire _2128;
    wire _2144;
    wire _2051;
    wire _2052;
    wire _2060;
    wire _2080;
    wire _2127;
    wire _2143;
    wire _2054;
    wire _2056;
    wire _2059;
    wire _2079;
    wire _2126;
    wire _2142;
    wire _2055;
    wire _2057;
    wire _2058;
    wire _2078;
    wire _2125;
    wire _2141;
    wire _2062;
    wire _2065;
    wire _2072;
    wire _2077;
    wire _2124;
    wire _2140;
    wire _2063;
    wire _2064;
    wire _2071;
    wire _2076;
    wire _2123;
    wire _2139;
    wire _2066;
    wire _2068;
    wire _2070;
    wire _2075;
    wire _2122;
    wire _2138;
    wire _2067;
    wire _2069;
    wire _2073;
    wire _2074;
    wire _2121;
    wire _2137;
    wire _2082;
    wire _2085;
    wire _2093;
    wire _2112;
    wire _2120;
    wire _2136;
    wire _2083;
    wire _2084;
    wire _2092;
    wire _2111;
    wire _2119;
    wire _2135;
    wire _2086;
    wire _2088;
    wire _2091;
    wire _2110;
    wire _2118;
    wire _2134;
    wire _2087;
    wire _2089;
    wire _2090;
    wire _2109;
    wire _2117;
    wire _2133;
    wire _2094;
    wire _2097;
    wire _2104;
    wire _2108;
    wire _2116;
    wire _2132;
    wire _2095;
    wire _2096;
    wire _2103;
    wire _2107;
    wire _2115;
    wire _2131;
    wire _2098;
    wire _2100;
    wire _2102;
    wire _2106;
    wire _2114;
    wire _2130;
    wire _1772;
    wire _1773;
    wire _2099;
    wire _1774;
    wire _2101;
    wire _1775;
    wire _2105;
    wire _1776;
    wire _2113;
    wire _1777;
    wire _2129;
    wire [63:0] _2161;
    wire _2162;
    wire _2163;
    wire [31:0] _2165 = 32'b00000000000000000000000000000000;
    wire gnd = 1'b0;
    wire [31:0] _2164 = 32'b00000000000000000000000000000000;
    reg [31:0] _2166;
    reg [31:0] _2343;

    /* logic */
    always @* begin
        case (ra2)
        0: _2342 <= _2166;
        1: _2342 <= _2171;
        2: _2342 <= _2176;
        3: _2342 <= _2181;
        4: _2342 <= _2186;
        5: _2342 <= _2191;
        6: _2342 <= _2196;
        7: _2342 <= _2201;
        8: _2342 <= _2206;
        9: _2342 <= _2211;
        10: _2342 <= _2216;
        11: _2342 <= _2221;
        12: _2342 <= _2226;
        13: _2342 <= _2231;
        14: _2342 <= _2236;
        15: _2342 <= _2241;
        16: _2342 <= _2246;
        17: _2342 <= _2251;
        18: _2342 <= _2256;
        19: _2342 <= _2261;
        20: _2342 <= _2266;
        21: _2342 <= _2271;
        22: _2342 <= _2276;
        23: _2342 <= _2281;
        24: _2342 <= _2286;
        25: _2342 <= _2291;
        26: _2342 <= _2296;
        27: _2342 <= _2301;
        28: _2342 <= _2306;
        29: _2342 <= _2311;
        30: _2342 <= _2316;
        31: _2342 <= _2321;
        32: _2342 <= _2326;
        33: _2342 <= _2331;
        34: _2342 <= _2336;
        default: _2342 <= _2341;
        endcase
    end
    assign _2337 = _2161[35:35];
    assign _2338 = wr & _2337;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2341 <= _2339;
        else
            if (_2338)
                _2341 <= d;
    end
    assign _2332 = _2161[34:34];
    assign _2333 = wr & _2332;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2336 <= _2334;
        else
            if (_2333)
                _2336 <= d;
    end
    assign _2327 = _2161[33:33];
    assign _2328 = wr & _2327;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2331 <= _2329;
        else
            if (_2328)
                _2331 <= d;
    end
    assign _2322 = _2161[32:32];
    assign _2323 = wr & _2322;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2326 <= _2324;
        else
            if (_2323)
                _2326 <= d;
    end
    assign _2317 = _2161[31:31];
    assign _2318 = wr & _2317;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2321 <= _2319;
        else
            if (_2318)
                _2321 <= d;
    end
    assign _2312 = _2161[30:30];
    assign _2313 = wr & _2312;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2316 <= _2314;
        else
            if (_2313)
                _2316 <= d;
    end
    assign _2307 = _2161[29:29];
    assign _2308 = wr & _2307;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2311 <= _2309;
        else
            if (_2308)
                _2311 <= d;
    end
    assign _2302 = _2161[28:28];
    assign _2303 = wr & _2302;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2306 <= _2304;
        else
            if (_2303)
                _2306 <= d;
    end
    assign _2297 = _2161[27:27];
    assign _2298 = wr & _2297;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2301 <= _2299;
        else
            if (_2298)
                _2301 <= d;
    end
    assign _2292 = _2161[26:26];
    assign _2293 = wr & _2292;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2296 <= _2294;
        else
            if (_2293)
                _2296 <= d;
    end
    assign _2287 = _2161[25:25];
    assign _2288 = wr & _2287;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2291 <= _2289;
        else
            if (_2288)
                _2291 <= d;
    end
    assign _2282 = _2161[24:24];
    assign _2283 = wr & _2282;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2286 <= _2284;
        else
            if (_2283)
                _2286 <= d;
    end
    assign _2277 = _2161[23:23];
    assign _2278 = wr & _2277;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2281 <= _2279;
        else
            if (_2278)
                _2281 <= d;
    end
    assign _2272 = _2161[22:22];
    assign _2273 = wr & _2272;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2276 <= _2274;
        else
            if (_2273)
                _2276 <= d;
    end
    assign _2267 = _2161[21:21];
    assign _2268 = wr & _2267;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2271 <= _2269;
        else
            if (_2268)
                _2271 <= d;
    end
    assign _2262 = _2161[20:20];
    assign _2263 = wr & _2262;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2266 <= _2264;
        else
            if (_2263)
                _2266 <= d;
    end
    assign _2257 = _2161[19:19];
    assign _2258 = wr & _2257;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2261 <= _2259;
        else
            if (_2258)
                _2261 <= d;
    end
    assign _2252 = _2161[18:18];
    assign _2253 = wr & _2252;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2256 <= _2254;
        else
            if (_2253)
                _2256 <= d;
    end
    assign _2247 = _2161[17:17];
    assign _2248 = wr & _2247;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2251 <= _2249;
        else
            if (_2248)
                _2251 <= d;
    end
    assign _2242 = _2161[16:16];
    assign _2243 = wr & _2242;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2246 <= _2244;
        else
            if (_2243)
                _2246 <= d;
    end
    assign _2237 = _2161[15:15];
    assign _2238 = wr & _2237;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2241 <= _2239;
        else
            if (_2238)
                _2241 <= d;
    end
    assign _2232 = _2161[14:14];
    assign _2233 = wr & _2232;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2236 <= _2234;
        else
            if (_2233)
                _2236 <= d;
    end
    assign _2227 = _2161[13:13];
    assign _2228 = wr & _2227;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2231 <= _2229;
        else
            if (_2228)
                _2231 <= d;
    end
    assign _2222 = _2161[12:12];
    assign _2223 = wr & _2222;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2226 <= _2224;
        else
            if (_2223)
                _2226 <= d;
    end
    assign _2217 = _2161[11:11];
    assign _2218 = wr & _2217;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2221 <= _2219;
        else
            if (_2218)
                _2221 <= d;
    end
    assign _2212 = _2161[10:10];
    assign _2213 = wr & _2212;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2216 <= _2214;
        else
            if (_2213)
                _2216 <= d;
    end
    assign _2207 = _2161[9:9];
    assign _2208 = wr & _2207;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2211 <= _2209;
        else
            if (_2208)
                _2211 <= d;
    end
    assign _2202 = _2161[8:8];
    assign _2203 = wr & _2202;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2206 <= _2204;
        else
            if (_2203)
                _2206 <= d;
    end
    assign _2197 = _2161[7:7];
    assign _2198 = wr & _2197;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2201 <= _2199;
        else
            if (_2198)
                _2201 <= d;
    end
    assign _2192 = _2161[6:6];
    assign _2193 = wr & _2192;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2196 <= _2194;
        else
            if (_2193)
                _2196 <= d;
    end
    assign _2187 = _2161[5:5];
    assign _2188 = wr & _2187;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2191 <= _2189;
        else
            if (_2188)
                _2191 <= d;
    end
    assign _2182 = _2161[4:4];
    assign _2183 = wr & _2182;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2186 <= _2184;
        else
            if (_2183)
                _2186 <= d;
    end
    assign _2177 = _2161[3:3];
    assign _2178 = wr & _2177;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2181 <= _2179;
        else
            if (_2178)
                _2181 <= d;
    end
    assign _2172 = _2161[2:2];
    assign _2173 = wr & _2172;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2176 <= _2174;
        else
            if (_2173)
                _2176 <= d;
    end
    assign _2167 = _2161[1:1];
    assign _2168 = wr & _2167;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2171 <= _2169;
        else
            if (_2168)
                _2171 <= d;
    end
    assign _1778 = ~ _1772;
    assign _1781 = _1779 & _1778;
    assign _1789 = _1785 & _1781;
    assign _1809 = _1801 & _1789;
    assign _1857 = _1841 & _1809;
    assign _1969 = _1937 & _1857;
    assign _1779 = ~ _1773;
    assign _1780 = _1779 & _1772;
    assign _1788 = _1785 & _1780;
    assign _1808 = _1801 & _1788;
    assign _1856 = _1841 & _1808;
    assign _1968 = _1937 & _1856;
    assign _1782 = ~ _1772;
    assign _1784 = _1773 & _1782;
    assign _1787 = _1785 & _1784;
    assign _1807 = _1801 & _1787;
    assign _1855 = _1841 & _1807;
    assign _1967 = _1937 & _1855;
    assign _1783 = _1773 & _1772;
    assign _1785 = ~ _1774;
    assign _1786 = _1785 & _1783;
    assign _1806 = _1801 & _1786;
    assign _1854 = _1841 & _1806;
    assign _1966 = _1937 & _1854;
    assign _1790 = ~ _1772;
    assign _1793 = _1791 & _1790;
    assign _1800 = _1774 & _1793;
    assign _1805 = _1801 & _1800;
    assign _1853 = _1841 & _1805;
    assign _1965 = _1937 & _1853;
    assign _1791 = ~ _1773;
    assign _1792 = _1791 & _1772;
    assign _1799 = _1774 & _1792;
    assign _1804 = _1801 & _1799;
    assign _1852 = _1841 & _1804;
    assign _1964 = _1937 & _1852;
    assign _1794 = ~ _1772;
    assign _1796 = _1773 & _1794;
    assign _1798 = _1774 & _1796;
    assign _1803 = _1801 & _1798;
    assign _1851 = _1841 & _1803;
    assign _1963 = _1937 & _1851;
    assign _1795 = _1773 & _1772;
    assign _1797 = _1774 & _1795;
    assign _1801 = ~ _1775;
    assign _1802 = _1801 & _1797;
    assign _1850 = _1841 & _1802;
    assign _1962 = _1937 & _1850;
    assign _1810 = ~ _1772;
    assign _1813 = _1811 & _1810;
    assign _1821 = _1817 & _1813;
    assign _1840 = _1775 & _1821;
    assign _1849 = _1841 & _1840;
    assign _1961 = _1937 & _1849;
    assign _1811 = ~ _1773;
    assign _1812 = _1811 & _1772;
    assign _1820 = _1817 & _1812;
    assign _1839 = _1775 & _1820;
    assign _1848 = _1841 & _1839;
    assign _1960 = _1937 & _1848;
    assign _1814 = ~ _1772;
    assign _1816 = _1773 & _1814;
    assign _1819 = _1817 & _1816;
    assign _1838 = _1775 & _1819;
    assign _1847 = _1841 & _1838;
    assign _1959 = _1937 & _1847;
    assign _1815 = _1773 & _1772;
    assign _1817 = ~ _1774;
    assign _1818 = _1817 & _1815;
    assign _1837 = _1775 & _1818;
    assign _1846 = _1841 & _1837;
    assign _1958 = _1937 & _1846;
    assign _1822 = ~ _1772;
    assign _1825 = _1823 & _1822;
    assign _1832 = _1774 & _1825;
    assign _1836 = _1775 & _1832;
    assign _1845 = _1841 & _1836;
    assign _1957 = _1937 & _1845;
    assign _1823 = ~ _1773;
    assign _1824 = _1823 & _1772;
    assign _1831 = _1774 & _1824;
    assign _1835 = _1775 & _1831;
    assign _1844 = _1841 & _1835;
    assign _1956 = _1937 & _1844;
    assign _1826 = ~ _1772;
    assign _1828 = _1773 & _1826;
    assign _1830 = _1774 & _1828;
    assign _1834 = _1775 & _1830;
    assign _1843 = _1841 & _1834;
    assign _1955 = _1937 & _1843;
    assign _1827 = _1773 & _1772;
    assign _1829 = _1774 & _1827;
    assign _1833 = _1775 & _1829;
    assign _1841 = ~ _1776;
    assign _1842 = _1841 & _1833;
    assign _1954 = _1937 & _1842;
    assign _1858 = ~ _1772;
    assign _1861 = _1859 & _1858;
    assign _1869 = _1865 & _1861;
    assign _1889 = _1881 & _1869;
    assign _1936 = _1776 & _1889;
    assign _1953 = _1937 & _1936;
    assign _1859 = ~ _1773;
    assign _1860 = _1859 & _1772;
    assign _1868 = _1865 & _1860;
    assign _1888 = _1881 & _1868;
    assign _1935 = _1776 & _1888;
    assign _1952 = _1937 & _1935;
    assign _1862 = ~ _1772;
    assign _1864 = _1773 & _1862;
    assign _1867 = _1865 & _1864;
    assign _1887 = _1881 & _1867;
    assign _1934 = _1776 & _1887;
    assign _1951 = _1937 & _1934;
    assign _1863 = _1773 & _1772;
    assign _1865 = ~ _1774;
    assign _1866 = _1865 & _1863;
    assign _1886 = _1881 & _1866;
    assign _1933 = _1776 & _1886;
    assign _1950 = _1937 & _1933;
    assign _1870 = ~ _1772;
    assign _1873 = _1871 & _1870;
    assign _1880 = _1774 & _1873;
    assign _1885 = _1881 & _1880;
    assign _1932 = _1776 & _1885;
    assign _1949 = _1937 & _1932;
    assign _1871 = ~ _1773;
    assign _1872 = _1871 & _1772;
    assign _1879 = _1774 & _1872;
    assign _1884 = _1881 & _1879;
    assign _1931 = _1776 & _1884;
    assign _1948 = _1937 & _1931;
    assign _1874 = ~ _1772;
    assign _1876 = _1773 & _1874;
    assign _1878 = _1774 & _1876;
    assign _1883 = _1881 & _1878;
    assign _1930 = _1776 & _1883;
    assign _1947 = _1937 & _1930;
    assign _1875 = _1773 & _1772;
    assign _1877 = _1774 & _1875;
    assign _1881 = ~ _1775;
    assign _1882 = _1881 & _1877;
    assign _1929 = _1776 & _1882;
    assign _1946 = _1937 & _1929;
    assign _1890 = ~ _1772;
    assign _1893 = _1891 & _1890;
    assign _1901 = _1897 & _1893;
    assign _1920 = _1775 & _1901;
    assign _1928 = _1776 & _1920;
    assign _1945 = _1937 & _1928;
    assign _1891 = ~ _1773;
    assign _1892 = _1891 & _1772;
    assign _1900 = _1897 & _1892;
    assign _1919 = _1775 & _1900;
    assign _1927 = _1776 & _1919;
    assign _1944 = _1937 & _1927;
    assign _1894 = ~ _1772;
    assign _1896 = _1773 & _1894;
    assign _1899 = _1897 & _1896;
    assign _1918 = _1775 & _1899;
    assign _1926 = _1776 & _1918;
    assign _1943 = _1937 & _1926;
    assign _1895 = _1773 & _1772;
    assign _1897 = ~ _1774;
    assign _1898 = _1897 & _1895;
    assign _1917 = _1775 & _1898;
    assign _1925 = _1776 & _1917;
    assign _1942 = _1937 & _1925;
    assign _1902 = ~ _1772;
    assign _1905 = _1903 & _1902;
    assign _1912 = _1774 & _1905;
    assign _1916 = _1775 & _1912;
    assign _1924 = _1776 & _1916;
    assign _1941 = _1937 & _1924;
    assign _1903 = ~ _1773;
    assign _1904 = _1903 & _1772;
    assign _1911 = _1774 & _1904;
    assign _1915 = _1775 & _1911;
    assign _1923 = _1776 & _1915;
    assign _1940 = _1937 & _1923;
    assign _1906 = ~ _1772;
    assign _1908 = _1773 & _1906;
    assign _1910 = _1774 & _1908;
    assign _1914 = _1775 & _1910;
    assign _1922 = _1776 & _1914;
    assign _1939 = _1937 & _1922;
    assign _1907 = _1773 & _1772;
    assign _1909 = _1774 & _1907;
    assign _1913 = _1775 & _1909;
    assign _1921 = _1776 & _1913;
    assign _1937 = ~ _1777;
    assign _1938 = _1937 & _1921;
    assign _1970 = ~ _1772;
    assign _1973 = _1971 & _1970;
    assign _1981 = _1977 & _1973;
    assign _2001 = _1993 & _1981;
    assign _2049 = _2033 & _2001;
    assign _2160 = _1777 & _2049;
    assign _1971 = ~ _1773;
    assign _1972 = _1971 & _1772;
    assign _1980 = _1977 & _1972;
    assign _2000 = _1993 & _1980;
    assign _2048 = _2033 & _2000;
    assign _2159 = _1777 & _2048;
    assign _1974 = ~ _1772;
    assign _1976 = _1773 & _1974;
    assign _1979 = _1977 & _1976;
    assign _1999 = _1993 & _1979;
    assign _2047 = _2033 & _1999;
    assign _2158 = _1777 & _2047;
    assign _1975 = _1773 & _1772;
    assign _1977 = ~ _1774;
    assign _1978 = _1977 & _1975;
    assign _1998 = _1993 & _1978;
    assign _2046 = _2033 & _1998;
    assign _2157 = _1777 & _2046;
    assign _1982 = ~ _1772;
    assign _1985 = _1983 & _1982;
    assign _1992 = _1774 & _1985;
    assign _1997 = _1993 & _1992;
    assign _2045 = _2033 & _1997;
    assign _2156 = _1777 & _2045;
    assign _1983 = ~ _1773;
    assign _1984 = _1983 & _1772;
    assign _1991 = _1774 & _1984;
    assign _1996 = _1993 & _1991;
    assign _2044 = _2033 & _1996;
    assign _2155 = _1777 & _2044;
    assign _1986 = ~ _1772;
    assign _1988 = _1773 & _1986;
    assign _1990 = _1774 & _1988;
    assign _1995 = _1993 & _1990;
    assign _2043 = _2033 & _1995;
    assign _2154 = _1777 & _2043;
    assign _1987 = _1773 & _1772;
    assign _1989 = _1774 & _1987;
    assign _1993 = ~ _1775;
    assign _1994 = _1993 & _1989;
    assign _2042 = _2033 & _1994;
    assign _2153 = _1777 & _2042;
    assign _2002 = ~ _1772;
    assign _2005 = _2003 & _2002;
    assign _2013 = _2009 & _2005;
    assign _2032 = _1775 & _2013;
    assign _2041 = _2033 & _2032;
    assign _2152 = _1777 & _2041;
    assign _2003 = ~ _1773;
    assign _2004 = _2003 & _1772;
    assign _2012 = _2009 & _2004;
    assign _2031 = _1775 & _2012;
    assign _2040 = _2033 & _2031;
    assign _2151 = _1777 & _2040;
    assign _2006 = ~ _1772;
    assign _2008 = _1773 & _2006;
    assign _2011 = _2009 & _2008;
    assign _2030 = _1775 & _2011;
    assign _2039 = _2033 & _2030;
    assign _2150 = _1777 & _2039;
    assign _2007 = _1773 & _1772;
    assign _2009 = ~ _1774;
    assign _2010 = _2009 & _2007;
    assign _2029 = _1775 & _2010;
    assign _2038 = _2033 & _2029;
    assign _2149 = _1777 & _2038;
    assign _2014 = ~ _1772;
    assign _2017 = _2015 & _2014;
    assign _2024 = _1774 & _2017;
    assign _2028 = _1775 & _2024;
    assign _2037 = _2033 & _2028;
    assign _2148 = _1777 & _2037;
    assign _2015 = ~ _1773;
    assign _2016 = _2015 & _1772;
    assign _2023 = _1774 & _2016;
    assign _2027 = _1775 & _2023;
    assign _2036 = _2033 & _2027;
    assign _2147 = _1777 & _2036;
    assign _2018 = ~ _1772;
    assign _2020 = _1773 & _2018;
    assign _2022 = _1774 & _2020;
    assign _2026 = _1775 & _2022;
    assign _2035 = _2033 & _2026;
    assign _2146 = _1777 & _2035;
    assign _2019 = _1773 & _1772;
    assign _2021 = _1774 & _2019;
    assign _2025 = _1775 & _2021;
    assign _2033 = ~ _1776;
    assign _2034 = _2033 & _2025;
    assign _2145 = _1777 & _2034;
    assign _2050 = ~ _1772;
    assign _2053 = _2051 & _2050;
    assign _2061 = _2057 & _2053;
    assign _2081 = _2073 & _2061;
    assign _2128 = _1776 & _2081;
    assign _2144 = _1777 & _2128;
    assign _2051 = ~ _1773;
    assign _2052 = _2051 & _1772;
    assign _2060 = _2057 & _2052;
    assign _2080 = _2073 & _2060;
    assign _2127 = _1776 & _2080;
    assign _2143 = _1777 & _2127;
    assign _2054 = ~ _1772;
    assign _2056 = _1773 & _2054;
    assign _2059 = _2057 & _2056;
    assign _2079 = _2073 & _2059;
    assign _2126 = _1776 & _2079;
    assign _2142 = _1777 & _2126;
    assign _2055 = _1773 & _1772;
    assign _2057 = ~ _1774;
    assign _2058 = _2057 & _2055;
    assign _2078 = _2073 & _2058;
    assign _2125 = _1776 & _2078;
    assign _2141 = _1777 & _2125;
    assign _2062 = ~ _1772;
    assign _2065 = _2063 & _2062;
    assign _2072 = _1774 & _2065;
    assign _2077 = _2073 & _2072;
    assign _2124 = _1776 & _2077;
    assign _2140 = _1777 & _2124;
    assign _2063 = ~ _1773;
    assign _2064 = _2063 & _1772;
    assign _2071 = _1774 & _2064;
    assign _2076 = _2073 & _2071;
    assign _2123 = _1776 & _2076;
    assign _2139 = _1777 & _2123;
    assign _2066 = ~ _1772;
    assign _2068 = _1773 & _2066;
    assign _2070 = _1774 & _2068;
    assign _2075 = _2073 & _2070;
    assign _2122 = _1776 & _2075;
    assign _2138 = _1777 & _2122;
    assign _2067 = _1773 & _1772;
    assign _2069 = _1774 & _2067;
    assign _2073 = ~ _1775;
    assign _2074 = _2073 & _2069;
    assign _2121 = _1776 & _2074;
    assign _2137 = _1777 & _2121;
    assign _2082 = ~ _1772;
    assign _2085 = _2083 & _2082;
    assign _2093 = _2089 & _2085;
    assign _2112 = _1775 & _2093;
    assign _2120 = _1776 & _2112;
    assign _2136 = _1777 & _2120;
    assign _2083 = ~ _1773;
    assign _2084 = _2083 & _1772;
    assign _2092 = _2089 & _2084;
    assign _2111 = _1775 & _2092;
    assign _2119 = _1776 & _2111;
    assign _2135 = _1777 & _2119;
    assign _2086 = ~ _1772;
    assign _2088 = _1773 & _2086;
    assign _2091 = _2089 & _2088;
    assign _2110 = _1775 & _2091;
    assign _2118 = _1776 & _2110;
    assign _2134 = _1777 & _2118;
    assign _2087 = _1773 & _1772;
    assign _2089 = ~ _1774;
    assign _2090 = _2089 & _2087;
    assign _2109 = _1775 & _2090;
    assign _2117 = _1776 & _2109;
    assign _2133 = _1777 & _2117;
    assign _2094 = ~ _1772;
    assign _2097 = _2095 & _2094;
    assign _2104 = _1774 & _2097;
    assign _2108 = _1775 & _2104;
    assign _2116 = _1776 & _2108;
    assign _2132 = _1777 & _2116;
    assign _2095 = ~ _1773;
    assign _2096 = _2095 & _1772;
    assign _2103 = _1774 & _2096;
    assign _2107 = _1775 & _2103;
    assign _2115 = _1776 & _2107;
    assign _2131 = _1777 & _2115;
    assign _2098 = ~ _1772;
    assign _2100 = _1773 & _2098;
    assign _2102 = _1774 & _2100;
    assign _2106 = _1775 & _2102;
    assign _2114 = _1776 & _2106;
    assign _2130 = _1777 & _2114;
    assign _1772 = wa[0:0];
    assign _1773 = wa[1:1];
    assign _2099 = _1773 & _1772;
    assign _1774 = wa[2:2];
    assign _2101 = _1774 & _2099;
    assign _1775 = wa[3:3];
    assign _2105 = _1775 & _2101;
    assign _1776 = wa[4:4];
    assign _2113 = _1776 & _2105;
    assign _1777 = wa[5:5];
    assign _2129 = _1777 & _2113;
    assign _2161 = { _2129, _2130, _2131, _2132, _2133, _2134, _2135, _2136, _2137, _2138, _2139, _2140, _2141, _2142, _2143, _2144, _2145, _2146, _2147, _2148, _2149, _2150, _2151, _2152, _2153, _2154, _2155, _2156, _2157, _2158, _2159, _2160, _1938, _1939, _1940, _1941, _1942, _1943, _1944, _1945, _1946, _1947, _1948, _1949, _1950, _1951, _1952, _1953, _1954, _1955, _1956, _1957, _1958, _1959, _1960, _1961, _1962, _1963, _1964, _1965, _1966, _1967, _1968, _1969 };
    assign _2162 = _2161[0:0];
    assign _2163 = wr & _2162;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2166 <= _2164;
        else
            if (_2163)
                _2166 <= d;
    end
    always @* begin
        case (ra1)
        0: _2343 <= _2166;
        1: _2343 <= _2171;
        2: _2343 <= _2176;
        3: _2343 <= _2181;
        4: _2343 <= _2186;
        5: _2343 <= _2191;
        6: _2343 <= _2196;
        7: _2343 <= _2201;
        8: _2343 <= _2206;
        9: _2343 <= _2211;
        10: _2343 <= _2216;
        11: _2343 <= _2221;
        12: _2343 <= _2226;
        13: _2343 <= _2231;
        14: _2343 <= _2236;
        15: _2343 <= _2241;
        16: _2343 <= _2246;
        17: _2343 <= _2251;
        18: _2343 <= _2256;
        19: _2343 <= _2261;
        20: _2343 <= _2266;
        21: _2343 <= _2271;
        22: _2343 <= _2276;
        23: _2343 <= _2281;
        24: _2343 <= _2286;
        25: _2343 <= _2291;
        26: _2343 <= _2296;
        27: _2343 <= _2301;
        28: _2343 <= _2306;
        29: _2343 <= _2311;
        30: _2343 <= _2316;
        31: _2343 <= _2321;
        32: _2343 <= _2326;
        33: _2343 <= _2331;
        34: _2343 <= _2336;
        default: _2343 <= _2341;
        endcase
    end

    /* aliases */

    /* output assignments */
    assign q1 = _2343;
    assign q2 = _2342;

endmodule
